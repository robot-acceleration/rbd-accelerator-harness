        bproc.minv_block_in_R1_C1_dqdPE1(minv[0][0]);
        bproc.minv_block_in_R2_C1_dqdPE1(minv[1][0]);
        bproc.minv_block_in_R3_C1_dqdPE1(minv[2][0]);
        bproc.minv_block_in_R4_C1_dqdPE1(minv[3][0]);
        bproc.minv_block_in_R5_C1_dqdPE1(minv[4][0]);
        bproc.minv_block_in_R6_C1_dqdPE1(minv[5][0]);
        bproc.minv_block_in_R7_C1_dqdPE1(minv[6][0]);

        bproc.minv_block_in_R1_C2_dqdPE1(minv[0][1]);
        bproc.minv_block_in_R2_C2_dqdPE1(minv[1][1]);
        bproc.minv_block_in_R3_C2_dqdPE1(minv[2][1]);
        bproc.minv_block_in_R4_C2_dqdPE1(minv[3][1]);
        bproc.minv_block_in_R5_C2_dqdPE1(minv[4][1]);
        bproc.minv_block_in_R6_C2_dqdPE1(minv[5][1]);
        bproc.minv_block_in_R7_C2_dqdPE1(minv[6][1]);

        bproc.minv_block_in_R1_C3_dqdPE1(minv[0][2]);
        bproc.minv_block_in_R2_C3_dqdPE1(minv[1][2]);
        bproc.minv_block_in_R3_C3_dqdPE1(minv[2][2]);
        bproc.minv_block_in_R4_C3_dqdPE1(minv[3][2]);
        bproc.minv_block_in_R5_C3_dqdPE1(minv[4][2]);
        bproc.minv_block_in_R6_C3_dqdPE1(minv[5][2]);
        bproc.minv_block_in_R7_C3_dqdPE1(minv[6][2]);

        bproc.minv_block_in_R1_C4_dqdPE1(minv[0][3]);
        bproc.minv_block_in_R2_C4_dqdPE1(minv[1][3]);
        bproc.minv_block_in_R3_C4_dqdPE1(minv[2][3]);
        bproc.minv_block_in_R4_C4_dqdPE1(minv[3][3]);
        bproc.minv_block_in_R5_C4_dqdPE1(minv[4][3]);
        bproc.minv_block_in_R6_C4_dqdPE1(minv[5][3]);
        bproc.minv_block_in_R7_C4_dqdPE1(minv[6][3]);

        bproc.minv_block_in_R1_C5_dqdPE1(minv[0][4]);
        bproc.minv_block_in_R2_C5_dqdPE1(minv[1][4]);
        bproc.minv_block_in_R3_C5_dqdPE1(minv[2][4]);
        bproc.minv_block_in_R4_C5_dqdPE1(minv[3][4]);
        bproc.minv_block_in_R5_C5_dqdPE1(minv[4][4]);
        bproc.minv_block_in_R6_C5_dqdPE1(minv[5][4]);
        bproc.minv_block_in_R7_C5_dqdPE1(minv[6][4]);

        bproc.minv_block_in_R1_C6_dqdPE1(minv[0][5]);
        bproc.minv_block_in_R2_C6_dqdPE1(minv[1][5]);
        bproc.minv_block_in_R3_C6_dqdPE1(minv[2][5]);
        bproc.minv_block_in_R4_C6_dqdPE1(minv[3][5]);
        bproc.minv_block_in_R5_C6_dqdPE1(minv[4][5]);
        bproc.minv_block_in_R6_C6_dqdPE1(minv[5][5]);
        bproc.minv_block_in_R7_C6_dqdPE1(minv[6][5]);

        bproc.minv_block_in_R1_C7_dqdPE1(minv[0][6]);
        bproc.minv_block_in_R2_C7_dqdPE1(minv[1][6]);
        bproc.minv_block_in_R3_C7_dqdPE1(minv[2][6]);
        bproc.minv_block_in_R4_C7_dqdPE1(minv[3][6]);
        bproc.minv_block_in_R5_C7_dqdPE1(minv[4][6]);
        bproc.minv_block_in_R6_C7_dqdPE1(minv[5][6]);
        bproc.minv_block_in_R7_C7_dqdPE1(minv[6][6]);

        bproc.dtau_vec_in_R1_dqdPE1(new_dtaudq[0][0]);
        bproc.dtau_vec_in_R2_dqdPE1(new_dtaudq[1][0]);
        bproc.dtau_vec_in_R3_dqdPE1(new_dtaudq[2][0]);
        bproc.dtau_vec_in_R4_dqdPE1(new_dtaudq[3][0]);
        bproc.dtau_vec_in_R5_dqdPE1(new_dtaudq[4][0]);
        bproc.dtau_vec_in_R6_dqdPE1(new_dtaudq[5][0]);
        bproc.dtau_vec_in_R7_dqdPE1(new_dtaudq[6][0]);

        bproc.minv_block_in_R1_C1_dqdPE2(minv[0][0]);
        bproc.minv_block_in_R2_C1_dqdPE2(minv[1][0]);
        bproc.minv_block_in_R3_C1_dqdPE2(minv[2][0]);
        bproc.minv_block_in_R4_C1_dqdPE2(minv[3][0]);
        bproc.minv_block_in_R5_C1_dqdPE2(minv[4][0]);
        bproc.minv_block_in_R6_C1_dqdPE2(minv[5][0]);
        bproc.minv_block_in_R7_C1_dqdPE2(minv[6][0]);

        bproc.minv_block_in_R1_C2_dqdPE2(minv[0][1]);
        bproc.minv_block_in_R2_C2_dqdPE2(minv[1][1]);
        bproc.minv_block_in_R3_C2_dqdPE2(minv[2][1]);
        bproc.minv_block_in_R4_C2_dqdPE2(minv[3][1]);
        bproc.minv_block_in_R5_C2_dqdPE2(minv[4][1]);
        bproc.minv_block_in_R6_C2_dqdPE2(minv[5][1]);
        bproc.minv_block_in_R7_C2_dqdPE2(minv[6][1]);

        bproc.minv_block_in_R1_C3_dqdPE2(minv[0][2]);
        bproc.minv_block_in_R2_C3_dqdPE2(minv[1][2]);
        bproc.minv_block_in_R3_C3_dqdPE2(minv[2][2]);
        bproc.minv_block_in_R4_C3_dqdPE2(minv[3][2]);
        bproc.minv_block_in_R5_C3_dqdPE2(minv[4][2]);
        bproc.minv_block_in_R6_C3_dqdPE2(minv[5][2]);
        bproc.minv_block_in_R7_C3_dqdPE2(minv[6][2]);

        bproc.minv_block_in_R1_C4_dqdPE2(minv[0][3]);
        bproc.minv_block_in_R2_C4_dqdPE2(minv[1][3]);
        bproc.minv_block_in_R3_C4_dqdPE2(minv[2][3]);
        bproc.minv_block_in_R4_C4_dqdPE2(minv[3][3]);
        bproc.minv_block_in_R5_C4_dqdPE2(minv[4][3]);
        bproc.minv_block_in_R6_C4_dqdPE2(minv[5][3]);
        bproc.minv_block_in_R7_C4_dqdPE2(minv[6][3]);

        bproc.minv_block_in_R1_C5_dqdPE2(minv[0][4]);
        bproc.minv_block_in_R2_C5_dqdPE2(minv[1][4]);
        bproc.minv_block_in_R3_C5_dqdPE2(minv[2][4]);
        bproc.minv_block_in_R4_C5_dqdPE2(minv[3][4]);
        bproc.minv_block_in_R5_C5_dqdPE2(minv[4][4]);
        bproc.minv_block_in_R6_C5_dqdPE2(minv[5][4]);
        bproc.minv_block_in_R7_C5_dqdPE2(minv[6][4]);

        bproc.minv_block_in_R1_C6_dqdPE2(minv[0][5]);
        bproc.minv_block_in_R2_C6_dqdPE2(minv[1][5]);
        bproc.minv_block_in_R3_C6_dqdPE2(minv[2][5]);
        bproc.minv_block_in_R4_C6_dqdPE2(minv[3][5]);
        bproc.minv_block_in_R5_C6_dqdPE2(minv[4][5]);
        bproc.minv_block_in_R6_C6_dqdPE2(minv[5][5]);
        bproc.minv_block_in_R7_C6_dqdPE2(minv[6][5]);

        bproc.minv_block_in_R1_C7_dqdPE2(minv[0][6]);
        bproc.minv_block_in_R2_C7_dqdPE2(minv[1][6]);
        bproc.minv_block_in_R3_C7_dqdPE2(minv[2][6]);
        bproc.minv_block_in_R4_C7_dqdPE2(minv[3][6]);
        bproc.minv_block_in_R5_C7_dqdPE2(minv[4][6]);
        bproc.minv_block_in_R6_C7_dqdPE2(minv[5][6]);
        bproc.minv_block_in_R7_C7_dqdPE2(minv[6][6]);

        bproc.dtau_vec_in_R1_dqdPE2(new_dtaudq[0][1]);
        bproc.dtau_vec_in_R2_dqdPE2(new_dtaudq[1][1]);
        bproc.dtau_vec_in_R3_dqdPE2(new_dtaudq[2][1]);
        bproc.dtau_vec_in_R4_dqdPE2(new_dtaudq[3][1]);
        bproc.dtau_vec_in_R5_dqdPE2(new_dtaudq[4][1]);
        bproc.dtau_vec_in_R6_dqdPE2(new_dtaudq[5][1]);
        bproc.dtau_vec_in_R7_dqdPE2(new_dtaudq[6][1]);

        bproc.minv_block_in_R1_C1_dqdPE3(minv[0][0]);
        bproc.minv_block_in_R2_C1_dqdPE3(minv[1][0]);
        bproc.minv_block_in_R3_C1_dqdPE3(minv[2][0]);
        bproc.minv_block_in_R4_C1_dqdPE3(minv[3][0]);
        bproc.minv_block_in_R5_C1_dqdPE3(minv[4][0]);
        bproc.minv_block_in_R6_C1_dqdPE3(minv[5][0]);
        bproc.minv_block_in_R7_C1_dqdPE3(minv[6][0]);

        bproc.minv_block_in_R1_C2_dqdPE3(minv[0][1]);
        bproc.minv_block_in_R2_C2_dqdPE3(minv[1][1]);
        bproc.minv_block_in_R3_C2_dqdPE3(minv[2][1]);
        bproc.minv_block_in_R4_C2_dqdPE3(minv[3][1]);
        bproc.minv_block_in_R5_C2_dqdPE3(minv[4][1]);
        bproc.minv_block_in_R6_C2_dqdPE3(minv[5][1]);
        bproc.minv_block_in_R7_C2_dqdPE3(minv[6][1]);

        bproc.minv_block_in_R1_C3_dqdPE3(minv[0][2]);
        bproc.minv_block_in_R2_C3_dqdPE3(minv[1][2]);
        bproc.minv_block_in_R3_C3_dqdPE3(minv[2][2]);
        bproc.minv_block_in_R4_C3_dqdPE3(minv[3][2]);
        bproc.minv_block_in_R5_C3_dqdPE3(minv[4][2]);
        bproc.minv_block_in_R6_C3_dqdPE3(minv[5][2]);
        bproc.minv_block_in_R7_C3_dqdPE3(minv[6][2]);

        bproc.minv_block_in_R1_C4_dqdPE3(minv[0][3]);
        bproc.minv_block_in_R2_C4_dqdPE3(minv[1][3]);
        bproc.minv_block_in_R3_C4_dqdPE3(minv[2][3]);
        bproc.minv_block_in_R4_C4_dqdPE3(minv[3][3]);
        bproc.minv_block_in_R5_C4_dqdPE3(minv[4][3]);
        bproc.minv_block_in_R6_C4_dqdPE3(minv[5][3]);
        bproc.minv_block_in_R7_C4_dqdPE3(minv[6][3]);

        bproc.minv_block_in_R1_C5_dqdPE3(minv[0][4]);
        bproc.minv_block_in_R2_C5_dqdPE3(minv[1][4]);
        bproc.minv_block_in_R3_C5_dqdPE3(minv[2][4]);
        bproc.minv_block_in_R4_C5_dqdPE3(minv[3][4]);
        bproc.minv_block_in_R5_C5_dqdPE3(minv[4][4]);
        bproc.minv_block_in_R6_C5_dqdPE3(minv[5][4]);
        bproc.minv_block_in_R7_C5_dqdPE3(minv[6][4]);

        bproc.minv_block_in_R1_C6_dqdPE3(minv[0][5]);
        bproc.minv_block_in_R2_C6_dqdPE3(minv[1][5]);
        bproc.minv_block_in_R3_C6_dqdPE3(minv[2][5]);
        bproc.minv_block_in_R4_C6_dqdPE3(minv[3][5]);
        bproc.minv_block_in_R5_C6_dqdPE3(minv[4][5]);
        bproc.minv_block_in_R6_C6_dqdPE3(minv[5][5]);
        bproc.minv_block_in_R7_C6_dqdPE3(minv[6][5]);

        bproc.minv_block_in_R1_C7_dqdPE3(minv[0][6]);
        bproc.minv_block_in_R2_C7_dqdPE3(minv[1][6]);
        bproc.minv_block_in_R3_C7_dqdPE3(minv[2][6]);
        bproc.minv_block_in_R4_C7_dqdPE3(minv[3][6]);
        bproc.minv_block_in_R5_C7_dqdPE3(minv[4][6]);
        bproc.minv_block_in_R6_C7_dqdPE3(minv[5][6]);
        bproc.minv_block_in_R7_C7_dqdPE3(minv[6][6]);

        bproc.dtau_vec_in_R1_dqdPE3(new_dtaudq[0][2]);
        bproc.dtau_vec_in_R2_dqdPE3(new_dtaudq[1][2]);
        bproc.dtau_vec_in_R3_dqdPE3(new_dtaudq[2][2]);
        bproc.dtau_vec_in_R4_dqdPE3(new_dtaudq[3][2]);
        bproc.dtau_vec_in_R5_dqdPE3(new_dtaudq[4][2]);
        bproc.dtau_vec_in_R6_dqdPE3(new_dtaudq[5][2]);
        bproc.dtau_vec_in_R7_dqdPE3(new_dtaudq[6][2]);

        bproc.minv_block_in_R1_C1_dqdPE4(minv[0][0]);
        bproc.minv_block_in_R2_C1_dqdPE4(minv[1][0]);
        bproc.minv_block_in_R3_C1_dqdPE4(minv[2][0]);
        bproc.minv_block_in_R4_C1_dqdPE4(minv[3][0]);
        bproc.minv_block_in_R5_C1_dqdPE4(minv[4][0]);
        bproc.minv_block_in_R6_C1_dqdPE4(minv[5][0]);
        bproc.minv_block_in_R7_C1_dqdPE4(minv[6][0]);

        bproc.minv_block_in_R1_C2_dqdPE4(minv[0][1]);
        bproc.minv_block_in_R2_C2_dqdPE4(minv[1][1]);
        bproc.minv_block_in_R3_C2_dqdPE4(minv[2][1]);
        bproc.minv_block_in_R4_C2_dqdPE4(minv[3][1]);
        bproc.minv_block_in_R5_C2_dqdPE4(minv[4][1]);
        bproc.minv_block_in_R6_C2_dqdPE4(minv[5][1]);
        bproc.minv_block_in_R7_C2_dqdPE4(minv[6][1]);

        bproc.minv_block_in_R1_C3_dqdPE4(minv[0][2]);
        bproc.minv_block_in_R2_C3_dqdPE4(minv[1][2]);
        bproc.minv_block_in_R3_C3_dqdPE4(minv[2][2]);
        bproc.minv_block_in_R4_C3_dqdPE4(minv[3][2]);
        bproc.minv_block_in_R5_C3_dqdPE4(minv[4][2]);
        bproc.minv_block_in_R6_C3_dqdPE4(minv[5][2]);
        bproc.minv_block_in_R7_C3_dqdPE4(minv[6][2]);

        bproc.minv_block_in_R1_C4_dqdPE4(minv[0][3]);
        bproc.minv_block_in_R2_C4_dqdPE4(minv[1][3]);
        bproc.minv_block_in_R3_C4_dqdPE4(minv[2][3]);
        bproc.minv_block_in_R4_C4_dqdPE4(minv[3][3]);
        bproc.minv_block_in_R5_C4_dqdPE4(minv[4][3]);
        bproc.minv_block_in_R6_C4_dqdPE4(minv[5][3]);
        bproc.minv_block_in_R7_C4_dqdPE4(minv[6][3]);

        bproc.minv_block_in_R1_C5_dqdPE4(minv[0][4]);
        bproc.minv_block_in_R2_C5_dqdPE4(minv[1][4]);
        bproc.minv_block_in_R3_C5_dqdPE4(minv[2][4]);
        bproc.minv_block_in_R4_C5_dqdPE4(minv[3][4]);
        bproc.minv_block_in_R5_C5_dqdPE4(minv[4][4]);
        bproc.minv_block_in_R6_C5_dqdPE4(minv[5][4]);
        bproc.minv_block_in_R7_C5_dqdPE4(minv[6][4]);

        bproc.minv_block_in_R1_C6_dqdPE4(minv[0][5]);
        bproc.minv_block_in_R2_C6_dqdPE4(minv[1][5]);
        bproc.minv_block_in_R3_C6_dqdPE4(minv[2][5]);
        bproc.minv_block_in_R4_C6_dqdPE4(minv[3][5]);
        bproc.minv_block_in_R5_C6_dqdPE4(minv[4][5]);
        bproc.minv_block_in_R6_C6_dqdPE4(minv[5][5]);
        bproc.minv_block_in_R7_C6_dqdPE4(minv[6][5]);

        bproc.minv_block_in_R1_C7_dqdPE4(minv[0][6]);
        bproc.minv_block_in_R2_C7_dqdPE4(minv[1][6]);
        bproc.minv_block_in_R3_C7_dqdPE4(minv[2][6]);
        bproc.minv_block_in_R4_C7_dqdPE4(minv[3][6]);
        bproc.minv_block_in_R5_C7_dqdPE4(minv[4][6]);
        bproc.minv_block_in_R6_C7_dqdPE4(minv[5][6]);
        bproc.minv_block_in_R7_C7_dqdPE4(minv[6][6]);

        bproc.dtau_vec_in_R1_dqdPE4(new_dtaudq[0][3]);
        bproc.dtau_vec_in_R2_dqdPE4(new_dtaudq[1][3]);
        bproc.dtau_vec_in_R3_dqdPE4(new_dtaudq[2][3]);
        bproc.dtau_vec_in_R4_dqdPE4(new_dtaudq[3][3]);
        bproc.dtau_vec_in_R5_dqdPE4(new_dtaudq[4][3]);
        bproc.dtau_vec_in_R6_dqdPE4(new_dtaudq[5][3]);
        bproc.dtau_vec_in_R7_dqdPE4(new_dtaudq[6][3]);

        bproc.minv_block_in_R1_C1_dqdPE5(minv[0][0]);
        bproc.minv_block_in_R2_C1_dqdPE5(minv[1][0]);
        bproc.minv_block_in_R3_C1_dqdPE5(minv[2][0]);
        bproc.minv_block_in_R4_C1_dqdPE5(minv[3][0]);
        bproc.minv_block_in_R5_C1_dqdPE5(minv[4][0]);
        bproc.minv_block_in_R6_C1_dqdPE5(minv[5][0]);
        bproc.minv_block_in_R7_C1_dqdPE5(minv[6][0]);

        bproc.minv_block_in_R1_C2_dqdPE5(minv[0][1]);
        bproc.minv_block_in_R2_C2_dqdPE5(minv[1][1]);
        bproc.minv_block_in_R3_C2_dqdPE5(minv[2][1]);
        bproc.minv_block_in_R4_C2_dqdPE5(minv[3][1]);
        bproc.minv_block_in_R5_C2_dqdPE5(minv[4][1]);
        bproc.minv_block_in_R6_C2_dqdPE5(minv[5][1]);
        bproc.minv_block_in_R7_C2_dqdPE5(minv[6][1]);

        bproc.minv_block_in_R1_C3_dqdPE5(minv[0][2]);
        bproc.minv_block_in_R2_C3_dqdPE5(minv[1][2]);
        bproc.minv_block_in_R3_C3_dqdPE5(minv[2][2]);
        bproc.minv_block_in_R4_C3_dqdPE5(minv[3][2]);
        bproc.minv_block_in_R5_C3_dqdPE5(minv[4][2]);
        bproc.minv_block_in_R6_C3_dqdPE5(minv[5][2]);
        bproc.minv_block_in_R7_C3_dqdPE5(minv[6][2]);

        bproc.minv_block_in_R1_C4_dqdPE5(minv[0][3]);
        bproc.minv_block_in_R2_C4_dqdPE5(minv[1][3]);
        bproc.minv_block_in_R3_C4_dqdPE5(minv[2][3]);
        bproc.minv_block_in_R4_C4_dqdPE5(minv[3][3]);
        bproc.minv_block_in_R5_C4_dqdPE5(minv[4][3]);
        bproc.minv_block_in_R6_C4_dqdPE5(minv[5][3]);
        bproc.minv_block_in_R7_C4_dqdPE5(minv[6][3]);

        bproc.minv_block_in_R1_C5_dqdPE5(minv[0][4]);
        bproc.minv_block_in_R2_C5_dqdPE5(minv[1][4]);
        bproc.minv_block_in_R3_C5_dqdPE5(minv[2][4]);
        bproc.minv_block_in_R4_C5_dqdPE5(minv[3][4]);
        bproc.minv_block_in_R5_C5_dqdPE5(minv[4][4]);
        bproc.minv_block_in_R6_C5_dqdPE5(minv[5][4]);
        bproc.minv_block_in_R7_C5_dqdPE5(minv[6][4]);

        bproc.minv_block_in_R1_C6_dqdPE5(minv[0][5]);
        bproc.minv_block_in_R2_C6_dqdPE5(minv[1][5]);
        bproc.minv_block_in_R3_C6_dqdPE5(minv[2][5]);
        bproc.minv_block_in_R4_C6_dqdPE5(minv[3][5]);
        bproc.minv_block_in_R5_C6_dqdPE5(minv[4][5]);
        bproc.minv_block_in_R6_C6_dqdPE5(minv[5][5]);
        bproc.minv_block_in_R7_C6_dqdPE5(minv[6][5]);

        bproc.minv_block_in_R1_C7_dqdPE5(minv[0][6]);
        bproc.minv_block_in_R2_C7_dqdPE5(minv[1][6]);
        bproc.minv_block_in_R3_C7_dqdPE5(minv[2][6]);
        bproc.minv_block_in_R4_C7_dqdPE5(minv[3][6]);
        bproc.minv_block_in_R5_C7_dqdPE5(minv[4][6]);
        bproc.minv_block_in_R6_C7_dqdPE5(minv[5][6]);
        bproc.minv_block_in_R7_C7_dqdPE5(minv[6][6]);

        bproc.dtau_vec_in_R1_dqdPE5(new_dtaudq[0][4]);
        bproc.dtau_vec_in_R2_dqdPE5(new_dtaudq[1][4]);
        bproc.dtau_vec_in_R3_dqdPE5(new_dtaudq[2][4]);
        bproc.dtau_vec_in_R4_dqdPE5(new_dtaudq[3][4]);
        bproc.dtau_vec_in_R5_dqdPE5(new_dtaudq[4][4]);
        bproc.dtau_vec_in_R6_dqdPE5(new_dtaudq[5][4]);
        bproc.dtau_vec_in_R7_dqdPE5(new_dtaudq[6][4]);

        bproc.minv_block_in_R1_C1_dqdPE6(minv[0][0]);
        bproc.minv_block_in_R2_C1_dqdPE6(minv[1][0]);
        bproc.minv_block_in_R3_C1_dqdPE6(minv[2][0]);
        bproc.minv_block_in_R4_C1_dqdPE6(minv[3][0]);
        bproc.minv_block_in_R5_C1_dqdPE6(minv[4][0]);
        bproc.minv_block_in_R6_C1_dqdPE6(minv[5][0]);
        bproc.minv_block_in_R7_C1_dqdPE6(minv[6][0]);

        bproc.minv_block_in_R1_C2_dqdPE6(minv[0][1]);
        bproc.minv_block_in_R2_C2_dqdPE6(minv[1][1]);
        bproc.minv_block_in_R3_C2_dqdPE6(minv[2][1]);
        bproc.minv_block_in_R4_C2_dqdPE6(minv[3][1]);
        bproc.minv_block_in_R5_C2_dqdPE6(minv[4][1]);
        bproc.minv_block_in_R6_C2_dqdPE6(minv[5][1]);
        bproc.minv_block_in_R7_C2_dqdPE6(minv[6][1]);

        bproc.minv_block_in_R1_C3_dqdPE6(minv[0][2]);
        bproc.minv_block_in_R2_C3_dqdPE6(minv[1][2]);
        bproc.minv_block_in_R3_C3_dqdPE6(minv[2][2]);
        bproc.minv_block_in_R4_C3_dqdPE6(minv[3][2]);
        bproc.minv_block_in_R5_C3_dqdPE6(minv[4][2]);
        bproc.minv_block_in_R6_C3_dqdPE6(minv[5][2]);
        bproc.minv_block_in_R7_C3_dqdPE6(minv[6][2]);

        bproc.minv_block_in_R1_C4_dqdPE6(minv[0][3]);
        bproc.minv_block_in_R2_C4_dqdPE6(minv[1][3]);
        bproc.minv_block_in_R3_C4_dqdPE6(minv[2][3]);
        bproc.minv_block_in_R4_C4_dqdPE6(minv[3][3]);
        bproc.minv_block_in_R5_C4_dqdPE6(minv[4][3]);
        bproc.minv_block_in_R6_C4_dqdPE6(minv[5][3]);
        bproc.minv_block_in_R7_C4_dqdPE6(minv[6][3]);

        bproc.minv_block_in_R1_C5_dqdPE6(minv[0][4]);
        bproc.minv_block_in_R2_C5_dqdPE6(minv[1][4]);
        bproc.minv_block_in_R3_C5_dqdPE6(minv[2][4]);
        bproc.minv_block_in_R4_C5_dqdPE6(minv[3][4]);
        bproc.minv_block_in_R5_C5_dqdPE6(minv[4][4]);
        bproc.minv_block_in_R6_C5_dqdPE6(minv[5][4]);
        bproc.minv_block_in_R7_C5_dqdPE6(minv[6][4]);

        bproc.minv_block_in_R1_C6_dqdPE6(minv[0][5]);
        bproc.minv_block_in_R2_C6_dqdPE6(minv[1][5]);
        bproc.minv_block_in_R3_C6_dqdPE6(minv[2][5]);
        bproc.minv_block_in_R4_C6_dqdPE6(minv[3][5]);
        bproc.minv_block_in_R5_C6_dqdPE6(minv[4][5]);
        bproc.minv_block_in_R6_C6_dqdPE6(minv[5][5]);
        bproc.minv_block_in_R7_C6_dqdPE6(minv[6][5]);

        bproc.minv_block_in_R1_C7_dqdPE6(minv[0][6]);
        bproc.minv_block_in_R2_C7_dqdPE6(minv[1][6]);
        bproc.minv_block_in_R3_C7_dqdPE6(minv[2][6]);
        bproc.minv_block_in_R4_C7_dqdPE6(minv[3][6]);
        bproc.minv_block_in_R5_C7_dqdPE6(minv[4][6]);
        bproc.minv_block_in_R6_C7_dqdPE6(minv[5][6]);
        bproc.minv_block_in_R7_C7_dqdPE6(minv[6][6]);

        bproc.dtau_vec_in_R1_dqdPE6(new_dtaudq[0][5]);
        bproc.dtau_vec_in_R2_dqdPE6(new_dtaudq[1][5]);
        bproc.dtau_vec_in_R3_dqdPE6(new_dtaudq[2][5]);
        bproc.dtau_vec_in_R4_dqdPE6(new_dtaudq[3][5]);
        bproc.dtau_vec_in_R5_dqdPE6(new_dtaudq[4][5]);
        bproc.dtau_vec_in_R6_dqdPE6(new_dtaudq[5][5]);
        bproc.dtau_vec_in_R7_dqdPE6(new_dtaudq[6][5]);

        bproc.minv_block_in_R1_C1_dqdPE7(minv[0][0]);
        bproc.minv_block_in_R2_C1_dqdPE7(minv[1][0]);
        bproc.minv_block_in_R3_C1_dqdPE7(minv[2][0]);
        bproc.minv_block_in_R4_C1_dqdPE7(minv[3][0]);
        bproc.minv_block_in_R5_C1_dqdPE7(minv[4][0]);
        bproc.minv_block_in_R6_C1_dqdPE7(minv[5][0]);
        bproc.minv_block_in_R7_C1_dqdPE7(minv[6][0]);

        bproc.minv_block_in_R1_C2_dqdPE7(minv[0][1]);
        bproc.minv_block_in_R2_C2_dqdPE7(minv[1][1]);
        bproc.minv_block_in_R3_C2_dqdPE7(minv[2][1]);
        bproc.minv_block_in_R4_C2_dqdPE7(minv[3][1]);
        bproc.minv_block_in_R5_C2_dqdPE7(minv[4][1]);
        bproc.minv_block_in_R6_C2_dqdPE7(minv[5][1]);
        bproc.minv_block_in_R7_C2_dqdPE7(minv[6][1]);

        bproc.minv_block_in_R1_C3_dqdPE7(minv[0][2]);
        bproc.minv_block_in_R2_C3_dqdPE7(minv[1][2]);
        bproc.minv_block_in_R3_C3_dqdPE7(minv[2][2]);
        bproc.minv_block_in_R4_C3_dqdPE7(minv[3][2]);
        bproc.minv_block_in_R5_C3_dqdPE7(minv[4][2]);
        bproc.minv_block_in_R6_C3_dqdPE7(minv[5][2]);
        bproc.minv_block_in_R7_C3_dqdPE7(minv[6][2]);

        bproc.minv_block_in_R1_C4_dqdPE7(minv[0][3]);
        bproc.minv_block_in_R2_C4_dqdPE7(minv[1][3]);
        bproc.minv_block_in_R3_C4_dqdPE7(minv[2][3]);
        bproc.minv_block_in_R4_C4_dqdPE7(minv[3][3]);
        bproc.minv_block_in_R5_C4_dqdPE7(minv[4][3]);
        bproc.minv_block_in_R6_C4_dqdPE7(minv[5][3]);
        bproc.minv_block_in_R7_C4_dqdPE7(minv[6][3]);

        bproc.minv_block_in_R1_C5_dqdPE7(minv[0][4]);
        bproc.minv_block_in_R2_C5_dqdPE7(minv[1][4]);
        bproc.minv_block_in_R3_C5_dqdPE7(minv[2][4]);
        bproc.minv_block_in_R4_C5_dqdPE7(minv[3][4]);
        bproc.minv_block_in_R5_C5_dqdPE7(minv[4][4]);
        bproc.minv_block_in_R6_C5_dqdPE7(minv[5][4]);
        bproc.minv_block_in_R7_C5_dqdPE7(minv[6][4]);

        bproc.minv_block_in_R1_C6_dqdPE7(minv[0][5]);
        bproc.minv_block_in_R2_C6_dqdPE7(minv[1][5]);
        bproc.minv_block_in_R3_C6_dqdPE7(minv[2][5]);
        bproc.minv_block_in_R4_C6_dqdPE7(minv[3][5]);
        bproc.minv_block_in_R5_C6_dqdPE7(minv[4][5]);
        bproc.minv_block_in_R6_C6_dqdPE7(minv[5][5]);
        bproc.minv_block_in_R7_C6_dqdPE7(minv[6][5]);

        bproc.minv_block_in_R1_C7_dqdPE7(minv[0][6]);
        bproc.minv_block_in_R2_C7_dqdPE7(minv[1][6]);
        bproc.minv_block_in_R3_C7_dqdPE7(minv[2][6]);
        bproc.minv_block_in_R4_C7_dqdPE7(minv[3][6]);
        bproc.minv_block_in_R5_C7_dqdPE7(minv[4][6]);
        bproc.minv_block_in_R6_C7_dqdPE7(minv[5][6]);
        bproc.minv_block_in_R7_C7_dqdPE7(minv[6][6]);

        bproc.dtau_vec_in_R1_dqdPE7(new_dtaudq[0][6]);
        bproc.dtau_vec_in_R2_dqdPE7(new_dtaudq[1][6]);
        bproc.dtau_vec_in_R3_dqdPE7(new_dtaudq[2][6]);
        bproc.dtau_vec_in_R4_dqdPE7(new_dtaudq[3][6]);
        bproc.dtau_vec_in_R5_dqdPE7(new_dtaudq[4][6]);
        bproc.dtau_vec_in_R6_dqdPE7(new_dtaudq[5][6]);
        bproc.dtau_vec_in_R7_dqdPE7(new_dtaudq[6][6]);

