if (idx_backward_feed == 0) begin
    link_in_curr_PE1 = 8;
    link_in_par_PE1 = 7;
    link_in_derv_PE1 = 1;
    link_in_curr_PE2 = 8;
    link_in_par_PE2 = 7;
    link_in_derv_PE2 = 2;
    link_in_curr_PE3 = 8;
    link_in_par_PE3 = 7;
    link_in_derv_PE3 = 3;
    link_in_curr_PE4 = 8;
    link_in_par_PE4 = 7;
    link_in_derv_PE4 = 4;
    link_in_curr_PE5 = 8;
    link_in_par_PE5 = 7;
    link_in_derv_PE5 = 5;
    link_in_curr_PE6 = 8;
    link_in_par_PE6 = 7;
    link_in_derv_PE6 = 6;
    link_in_curr_PE7 = 8;
    link_in_par_PE7 = 7;
    link_in_derv_PE7 = 7;
end
else if (idx_backward_feed == 1) begin
    link_in_curr_PE1 = 7;
    link_in_par_PE1 = 6;
    link_in_derv_PE1 = 1;
    link_in_curr_PE2 = 7;
    link_in_par_PE2 = 6;
    link_in_derv_PE2 = 2;
    link_in_curr_PE3 = 7;
    link_in_par_PE3 = 6;
    link_in_derv_PE3 = 3;
    link_in_curr_PE4 = 7;
    link_in_par_PE4 = 6;
    link_in_derv_PE4 = 4;
    link_in_curr_PE5 = 7;
    link_in_par_PE5 = 6;
    link_in_derv_PE5 = 5;
    link_in_curr_PE6 = 7;
    link_in_par_PE6 = 6;
    link_in_derv_PE6 = 6;
    link_in_curr_PE7 = 7;
    link_in_par_PE7 = 6;
    link_in_derv_PE7 = 7;
end
else if (idx_backward_feed == 2) begin
    link_in_curr_PE1 = 6;
    link_in_par_PE1 = 5;
    link_in_derv_PE1 = 1;
    link_in_curr_PE2 = 6;
    link_in_par_PE2 = 5;
    link_in_derv_PE2 = 2;
    link_in_curr_PE3 = 6;
    link_in_par_PE3 = 5;
    link_in_derv_PE3 = 3;
    link_in_curr_PE4 = 6;
    link_in_par_PE4 = 5;
    link_in_derv_PE4 = 4;
    link_in_curr_PE5 = 6;
    link_in_par_PE5 = 5;
    link_in_derv_PE5 = 5;
    link_in_curr_PE6 = 6;
    link_in_par_PE6 = 5;
    link_in_derv_PE6 = 6;
    link_in_curr_PE7 = 6;
    link_in_par_PE7 = 5;
    link_in_derv_PE7 = 7;
end
else if (idx_backward_feed == 3) begin
    link_in_curr_PE1 = 5;
    link_in_par_PE1 = 4;
    link_in_derv_PE1 = 1;
    link_in_curr_PE2 = 5;
    link_in_par_PE2 = 4;
    link_in_derv_PE2 = 2;
    link_in_curr_PE3 = 5;
    link_in_par_PE3 = 4;
    link_in_derv_PE3 = 3;
    link_in_curr_PE4 = 5;
    link_in_par_PE4 = 4;
    link_in_derv_PE4 = 4;
    link_in_curr_PE5 = 5;
    link_in_par_PE5 = 4;
    link_in_derv_PE5 = 5;
    link_in_curr_PE6 = 5;
    link_in_par_PE6 = 4;
    link_in_derv_PE6 = 6;
    link_in_curr_PE7 = 5;
    link_in_par_PE7 = 4;
    link_in_derv_PE7 = 7;
end
else if (idx_backward_feed == 4) begin
    link_in_curr_PE1 = 4;
    link_in_par_PE1 = 3;
    link_in_derv_PE1 = 1;
    link_in_curr_PE2 = 4;
    link_in_par_PE2 = 3;
    link_in_derv_PE2 = 2;
    link_in_curr_PE3 = 4;
    link_in_par_PE3 = 3;
    link_in_derv_PE3 = 3;
    link_in_curr_PE4 = 4;
    link_in_par_PE4 = 3;
    link_in_derv_PE4 = 4;
    link_in_curr_PE5 = 4;
    link_in_par_PE5 = 3;
    link_in_derv_PE5 = 5;
    link_in_curr_PE6 = 4;
    link_in_par_PE6 = 3;
    link_in_derv_PE6 = 6;
    link_in_curr_PE7 = 4;
    link_in_par_PE7 = 3;
    link_in_derv_PE7 = 7;
end
else if (idx_backward_feed == 5) begin
    link_in_curr_PE1 = 3;
    link_in_par_PE1 = 2;
    link_in_derv_PE1 = 1;
    link_in_curr_PE2 = 3;
    link_in_par_PE2 = 2;
    link_in_derv_PE2 = 2;
    link_in_curr_PE3 = 3;
    link_in_par_PE3 = 2;
    link_in_derv_PE3 = 3;
    link_in_curr_PE4 = 3;
    link_in_par_PE4 = 2;
    link_in_derv_PE4 = 4;
    link_in_curr_PE5 = 3;
    link_in_par_PE5 = 2;
    link_in_derv_PE5 = 5;
    link_in_curr_PE6 = 3;
    link_in_par_PE6 = 2;
    link_in_derv_PE6 = 6;
    link_in_curr_PE7 = 3;
    link_in_par_PE7 = 2;
    link_in_derv_PE7 = 7;
end
else if (idx_backward_feed == 6) begin
    link_in_curr_PE1 = 2;
    link_in_par_PE1 = 1;
    link_in_derv_PE1 = 1;
    link_in_curr_PE2 = 2;
    link_in_par_PE2 = 1;
    link_in_derv_PE2 = 2;
    link_in_curr_PE3 = 2;
    link_in_par_PE3 = 1;
    link_in_derv_PE3 = 3;
    link_in_curr_PE4 = 2;
    link_in_par_PE4 = 1;
    link_in_derv_PE4 = 4;
    link_in_curr_PE5 = 2;
    link_in_par_PE5 = 1;
    link_in_derv_PE5 = 5;
    link_in_curr_PE6 = 2;
    link_in_par_PE6 = 1;
    link_in_derv_PE6 = 6;
    link_in_curr_PE7 = 2;
    link_in_par_PE7 = 1;
    link_in_derv_PE7 = 7;
end
else if (idx_backward_feed == 7) begin
    link_in_curr_PE1 = 1;
    link_in_par_PE1 = 0;
    link_in_derv_PE1 = 1;
    link_in_curr_PE2 = 1;
    link_in_par_PE2 = 0;
    link_in_derv_PE2 = 2;
    link_in_curr_PE3 = 1;
    link_in_par_PE3 = 0;
    link_in_derv_PE3 = 3;
    link_in_curr_PE4 = 1;
    link_in_par_PE4 = 0;
    link_in_derv_PE4 = 4;
    link_in_curr_PE5 = 1;
    link_in_par_PE5 = 0;
    link_in_derv_PE5 = 5;
    link_in_curr_PE6 = 1;
    link_in_par_PE6 = 0;
    link_in_derv_PE6 = 6;
    link_in_curr_PE7 = 1;
    link_in_par_PE7 = 0;
    link_in_derv_PE7 = 7;
end
