import Clocks::*;
(* always_ready, always_enabled *)
interface FProc;
    (* always_ready *)
    method Action get_data();

    //-------- RNEA INPUTS -----

    method Action link_in_rnea(Bit#(3) v);
    method Action sinq_val_in_rnea(Bit#(32) v);
    method Action cosq_val_in_rnea(Bit#(32) v);

    method Action qd_val_in_rnea(Bit#(32) v);
    method Action qdd_val_in_rnea(Bit#(32) v);

    method Action v_prev_vec_in_AX_rnea(Bit#(32) v);
    method Action v_prev_vec_in_AY_rnea(Bit#(32) v);
    method Action v_prev_vec_in_AZ_rnea(Bit#(32) v);
    method Action v_prev_vec_in_LX_rnea(Bit#(32) v);
    method Action v_prev_vec_in_LY_rnea(Bit#(32) v);
    method Action v_prev_vec_in_LZ_rnea(Bit#(32) v);
    method Action a_prev_vec_in_AX_rnea(Bit#(32) v);
    method Action a_prev_vec_in_AY_rnea(Bit#(32) v);
    method Action a_prev_vec_in_AZ_rnea(Bit#(32) v);
    method Action a_prev_vec_in_LX_rnea(Bit#(32) v);
    method Action a_prev_vec_in_LY_rnea(Bit#(32) v);
    method Action a_prev_vec_in_LZ_rnea(Bit#(32) v);

   //--------------------------

    //-------- DQ AND DQD INPUTS -----

    method Action link_in_dqPE1(Bit#(3) v);
    method Action link_in_dqPE2(Bit#(3) v);
    method Action link_in_dqPE3(Bit#(3) v);
    method Action link_in_dqPE4(Bit#(3) v);
    method Action link_in_dqPE5(Bit#(3) v);
    method Action link_in_dqPE6(Bit#(3) v);
    method Action link_in_dqPE7(Bit#(3) v);
    method Action link_in_dqdPE1(Bit#(3) v);
    method Action link_in_dqdPE2(Bit#(3) v);
    method Action link_in_dqdPE3(Bit#(3) v);
    method Action link_in_dqdPE4(Bit#(3) v);
    method Action link_in_dqdPE5(Bit#(3) v);
    method Action link_in_dqdPE6(Bit#(3) v);
    method Action link_in_dqdPE7(Bit#(3) v);
    method Action derv_in_dqPE1(Bit#(3) v);
    method Action derv_in_dqPE2(Bit#(3) v);
    method Action derv_in_dqPE3(Bit#(3) v);
    method Action derv_in_dqPE4(Bit#(3) v);
    method Action derv_in_dqPE5(Bit#(3) v);
    method Action derv_in_dqPE6(Bit#(3) v);
    method Action derv_in_dqPE7(Bit#(3) v);
    method Action derv_in_dqdPE1(Bit#(3) v);
    method Action derv_in_dqdPE2(Bit#(3) v);
    method Action derv_in_dqdPE3(Bit#(3) v);
    method Action derv_in_dqdPE4(Bit#(3) v);
    method Action derv_in_dqdPE5(Bit#(3) v);
    method Action derv_in_dqdPE6(Bit#(3) v);
    method Action derv_in_dqdPE7(Bit#(3) v);

    method Action sinq_val_in_dqPE1(Bit#(32) v);
    method Action sinq_val_in_dqPE2(Bit#(32) v);
    method Action sinq_val_in_dqPE3(Bit#(32) v);
    method Action sinq_val_in_dqPE4(Bit#(32) v);
    method Action sinq_val_in_dqPE5(Bit#(32) v);
    method Action sinq_val_in_dqPE6(Bit#(32) v);
    method Action sinq_val_in_dqPE7(Bit#(32) v);
    method Action sinq_val_in_dqdPE1(Bit#(32) v);
    method Action sinq_val_in_dqdPE2(Bit#(32) v);
    method Action sinq_val_in_dqdPE3(Bit#(32) v);
    method Action sinq_val_in_dqdPE4(Bit#(32) v);
    method Action sinq_val_in_dqdPE5(Bit#(32) v);
    method Action sinq_val_in_dqdPE6(Bit#(32) v);
    method Action sinq_val_in_dqdPE7(Bit#(32) v);
    method Action cosq_val_in_dqPE1(Bit#(32) v);
    method Action cosq_val_in_dqPE2(Bit#(32) v);
    method Action cosq_val_in_dqPE3(Bit#(32) v);
    method Action cosq_val_in_dqPE4(Bit#(32) v);
    method Action cosq_val_in_dqPE5(Bit#(32) v);
    method Action cosq_val_in_dqPE6(Bit#(32) v);
    method Action cosq_val_in_dqPE7(Bit#(32) v);
    method Action cosq_val_in_dqdPE1(Bit#(32) v);
    method Action cosq_val_in_dqdPE2(Bit#(32) v);
    method Action cosq_val_in_dqdPE3(Bit#(32) v);
    method Action cosq_val_in_dqdPE4(Bit#(32) v);
    method Action cosq_val_in_dqdPE5(Bit#(32) v);
    method Action cosq_val_in_dqdPE6(Bit#(32) v);
    method Action cosq_val_in_dqdPE7(Bit#(32) v);
    method Action qd_val_in_dqPE1(Bit#(32) v);
    method Action qd_val_in_dqPE2(Bit#(32) v);
    method Action qd_val_in_dqPE3(Bit#(32) v);
    method Action qd_val_in_dqPE4(Bit#(32) v);
    method Action qd_val_in_dqPE5(Bit#(32) v);
    method Action qd_val_in_dqPE6(Bit#(32) v);
    method Action qd_val_in_dqPE7(Bit#(32) v);
    method Action qd_val_in_dqdPE1(Bit#(32) v);
    method Action qd_val_in_dqdPE2(Bit#(32) v);
    method Action qd_val_in_dqdPE3(Bit#(32) v);
    method Action qd_val_in_dqdPE4(Bit#(32) v);
    method Action qd_val_in_dqdPE5(Bit#(32) v);
    method Action qd_val_in_dqdPE6(Bit#(32) v);
    method Action qd_val_in_dqdPE7(Bit#(32) v);

    method Action v_curr_vec_in_AX_dqPE1(Bit#(32) v);
    method Action v_curr_vec_in_AY_dqPE1(Bit#(32) v);
    method Action v_curr_vec_in_AZ_dqPE1(Bit#(32) v);
    method Action v_curr_vec_in_LX_dqPE1(Bit#(32) v);
    method Action v_curr_vec_in_LY_dqPE1(Bit#(32) v);
    method Action v_curr_vec_in_LZ_dqPE1(Bit#(32) v);
    method Action v_curr_vec_in_AX_dqPE2(Bit#(32) v);
    method Action v_curr_vec_in_AY_dqPE2(Bit#(32) v);
    method Action v_curr_vec_in_AZ_dqPE2(Bit#(32) v);
    method Action v_curr_vec_in_LX_dqPE2(Bit#(32) v);
    method Action v_curr_vec_in_LY_dqPE2(Bit#(32) v);
    method Action v_curr_vec_in_LZ_dqPE2(Bit#(32) v);
    method Action v_curr_vec_in_AX_dqPE3(Bit#(32) v);
    method Action v_curr_vec_in_AY_dqPE3(Bit#(32) v);
    method Action v_curr_vec_in_AZ_dqPE3(Bit#(32) v);
    method Action v_curr_vec_in_LX_dqPE3(Bit#(32) v);
    method Action v_curr_vec_in_LY_dqPE3(Bit#(32) v);
    method Action v_curr_vec_in_LZ_dqPE3(Bit#(32) v);
    method Action v_curr_vec_in_AX_dqPE4(Bit#(32) v);
    method Action v_curr_vec_in_AY_dqPE4(Bit#(32) v);
    method Action v_curr_vec_in_AZ_dqPE4(Bit#(32) v);
    method Action v_curr_vec_in_LX_dqPE4(Bit#(32) v);
    method Action v_curr_vec_in_LY_dqPE4(Bit#(32) v);
    method Action v_curr_vec_in_LZ_dqPE4(Bit#(32) v);
    method Action v_curr_vec_in_AX_dqPE5(Bit#(32) v);
    method Action v_curr_vec_in_AY_dqPE5(Bit#(32) v);
    method Action v_curr_vec_in_AZ_dqPE5(Bit#(32) v);
    method Action v_curr_vec_in_LX_dqPE5(Bit#(32) v);
    method Action v_curr_vec_in_LY_dqPE5(Bit#(32) v);
    method Action v_curr_vec_in_LZ_dqPE5(Bit#(32) v);
    method Action v_curr_vec_in_AX_dqPE6(Bit#(32) v);
    method Action v_curr_vec_in_AY_dqPE6(Bit#(32) v);
    method Action v_curr_vec_in_AZ_dqPE6(Bit#(32) v);
    method Action v_curr_vec_in_LX_dqPE6(Bit#(32) v);
    method Action v_curr_vec_in_LY_dqPE6(Bit#(32) v);
    method Action v_curr_vec_in_LZ_dqPE6(Bit#(32) v);
    method Action v_curr_vec_in_AX_dqPE7(Bit#(32) v);
    method Action v_curr_vec_in_AY_dqPE7(Bit#(32) v);
    method Action v_curr_vec_in_AZ_dqPE7(Bit#(32) v);
    method Action v_curr_vec_in_LX_dqPE7(Bit#(32) v);
    method Action v_curr_vec_in_LY_dqPE7(Bit#(32) v);
    method Action v_curr_vec_in_LZ_dqPE7(Bit#(32) v);
    method Action v_curr_vec_in_AX_dqdPE1(Bit#(32) v);
    method Action v_curr_vec_in_AY_dqdPE1(Bit#(32) v);
    method Action v_curr_vec_in_AZ_dqdPE1(Bit#(32) v);
    method Action v_curr_vec_in_LX_dqdPE1(Bit#(32) v);
    method Action v_curr_vec_in_LY_dqdPE1(Bit#(32) v);
    method Action v_curr_vec_in_LZ_dqdPE1(Bit#(32) v);
    method Action v_curr_vec_in_AX_dqdPE2(Bit#(32) v);
    method Action v_curr_vec_in_AY_dqdPE2(Bit#(32) v);
    method Action v_curr_vec_in_AZ_dqdPE2(Bit#(32) v);
    method Action v_curr_vec_in_LX_dqdPE2(Bit#(32) v);
    method Action v_curr_vec_in_LY_dqdPE2(Bit#(32) v);
    method Action v_curr_vec_in_LZ_dqdPE2(Bit#(32) v);
    method Action v_curr_vec_in_AX_dqdPE3(Bit#(32) v);
    method Action v_curr_vec_in_AY_dqdPE3(Bit#(32) v);
    method Action v_curr_vec_in_AZ_dqdPE3(Bit#(32) v);
    method Action v_curr_vec_in_LX_dqdPE3(Bit#(32) v);
    method Action v_curr_vec_in_LY_dqdPE3(Bit#(32) v);
    method Action v_curr_vec_in_LZ_dqdPE3(Bit#(32) v);
    method Action v_curr_vec_in_AX_dqdPE4(Bit#(32) v);
    method Action v_curr_vec_in_AY_dqdPE4(Bit#(32) v);
    method Action v_curr_vec_in_AZ_dqdPE4(Bit#(32) v);
    method Action v_curr_vec_in_LX_dqdPE4(Bit#(32) v);
    method Action v_curr_vec_in_LY_dqdPE4(Bit#(32) v);
    method Action v_curr_vec_in_LZ_dqdPE4(Bit#(32) v);
    method Action v_curr_vec_in_AX_dqdPE5(Bit#(32) v);
    method Action v_curr_vec_in_AY_dqdPE5(Bit#(32) v);
    method Action v_curr_vec_in_AZ_dqdPE5(Bit#(32) v);
    method Action v_curr_vec_in_LX_dqdPE5(Bit#(32) v);
    method Action v_curr_vec_in_LY_dqdPE5(Bit#(32) v);
    method Action v_curr_vec_in_LZ_dqdPE5(Bit#(32) v);
    method Action v_curr_vec_in_AX_dqdPE6(Bit#(32) v);
    method Action v_curr_vec_in_AY_dqdPE6(Bit#(32) v);
    method Action v_curr_vec_in_AZ_dqdPE6(Bit#(32) v);
    method Action v_curr_vec_in_LX_dqdPE6(Bit#(32) v);
    method Action v_curr_vec_in_LY_dqdPE6(Bit#(32) v);
    method Action v_curr_vec_in_LZ_dqdPE6(Bit#(32) v);
    method Action v_curr_vec_in_AX_dqdPE7(Bit#(32) v);
    method Action v_curr_vec_in_AY_dqdPE7(Bit#(32) v);
    method Action v_curr_vec_in_AZ_dqdPE7(Bit#(32) v);
    method Action v_curr_vec_in_LX_dqdPE7(Bit#(32) v);
    method Action v_curr_vec_in_LY_dqdPE7(Bit#(32) v);
    method Action v_curr_vec_in_LZ_dqdPE7(Bit#(32) v);
    method Action a_curr_vec_in_AX_dqPE1(Bit#(32) v);
    method Action a_curr_vec_in_AY_dqPE1(Bit#(32) v);
    method Action a_curr_vec_in_AZ_dqPE1(Bit#(32) v);
    method Action a_curr_vec_in_LX_dqPE1(Bit#(32) v);
    method Action a_curr_vec_in_LY_dqPE1(Bit#(32) v);
    method Action a_curr_vec_in_LZ_dqPE1(Bit#(32) v);
    method Action a_curr_vec_in_AX_dqPE2(Bit#(32) v);
    method Action a_curr_vec_in_AY_dqPE2(Bit#(32) v);
    method Action a_curr_vec_in_AZ_dqPE2(Bit#(32) v);
    method Action a_curr_vec_in_LX_dqPE2(Bit#(32) v);
    method Action a_curr_vec_in_LY_dqPE2(Bit#(32) v);
    method Action a_curr_vec_in_LZ_dqPE2(Bit#(32) v);
    method Action a_curr_vec_in_AX_dqPE3(Bit#(32) v);
    method Action a_curr_vec_in_AY_dqPE3(Bit#(32) v);
    method Action a_curr_vec_in_AZ_dqPE3(Bit#(32) v);
    method Action a_curr_vec_in_LX_dqPE3(Bit#(32) v);
    method Action a_curr_vec_in_LY_dqPE3(Bit#(32) v);
    method Action a_curr_vec_in_LZ_dqPE3(Bit#(32) v);
    method Action a_curr_vec_in_AX_dqPE4(Bit#(32) v);
    method Action a_curr_vec_in_AY_dqPE4(Bit#(32) v);
    method Action a_curr_vec_in_AZ_dqPE4(Bit#(32) v);
    method Action a_curr_vec_in_LX_dqPE4(Bit#(32) v);
    method Action a_curr_vec_in_LY_dqPE4(Bit#(32) v);
    method Action a_curr_vec_in_LZ_dqPE4(Bit#(32) v);
    method Action a_curr_vec_in_AX_dqPE5(Bit#(32) v);
    method Action a_curr_vec_in_AY_dqPE5(Bit#(32) v);
    method Action a_curr_vec_in_AZ_dqPE5(Bit#(32) v);
    method Action a_curr_vec_in_LX_dqPE5(Bit#(32) v);
    method Action a_curr_vec_in_LY_dqPE5(Bit#(32) v);
    method Action a_curr_vec_in_LZ_dqPE5(Bit#(32) v);
    method Action a_curr_vec_in_AX_dqPE6(Bit#(32) v);
    method Action a_curr_vec_in_AY_dqPE6(Bit#(32) v);
    method Action a_curr_vec_in_AZ_dqPE6(Bit#(32) v);
    method Action a_curr_vec_in_LX_dqPE6(Bit#(32) v);
    method Action a_curr_vec_in_LY_dqPE6(Bit#(32) v);
    method Action a_curr_vec_in_LZ_dqPE6(Bit#(32) v);
    method Action a_curr_vec_in_AX_dqPE7(Bit#(32) v);
    method Action a_curr_vec_in_AY_dqPE7(Bit#(32) v);
    method Action a_curr_vec_in_AZ_dqPE7(Bit#(32) v);
    method Action a_curr_vec_in_LX_dqPE7(Bit#(32) v);
    method Action a_curr_vec_in_LY_dqPE7(Bit#(32) v);
    method Action a_curr_vec_in_LZ_dqPE7(Bit#(32) v);
    method Action a_curr_vec_in_AX_dqdPE1(Bit#(32) v);
    method Action a_curr_vec_in_AY_dqdPE1(Bit#(32) v);
    method Action a_curr_vec_in_AZ_dqdPE1(Bit#(32) v);
    method Action a_curr_vec_in_LX_dqdPE1(Bit#(32) v);
    method Action a_curr_vec_in_LY_dqdPE1(Bit#(32) v);
    method Action a_curr_vec_in_LZ_dqdPE1(Bit#(32) v);
    method Action a_curr_vec_in_AX_dqdPE2(Bit#(32) v);
    method Action a_curr_vec_in_AY_dqdPE2(Bit#(32) v);
    method Action a_curr_vec_in_AZ_dqdPE2(Bit#(32) v);
    method Action a_curr_vec_in_LX_dqdPE2(Bit#(32) v);
    method Action a_curr_vec_in_LY_dqdPE2(Bit#(32) v);
    method Action a_curr_vec_in_LZ_dqdPE2(Bit#(32) v);
    method Action a_curr_vec_in_AX_dqdPE3(Bit#(32) v);
    method Action a_curr_vec_in_AY_dqdPE3(Bit#(32) v);
    method Action a_curr_vec_in_AZ_dqdPE3(Bit#(32) v);
    method Action a_curr_vec_in_LX_dqdPE3(Bit#(32) v);
    method Action a_curr_vec_in_LY_dqdPE3(Bit#(32) v);
    method Action a_curr_vec_in_LZ_dqdPE3(Bit#(32) v);
    method Action a_curr_vec_in_AX_dqdPE4(Bit#(32) v);
    method Action a_curr_vec_in_AY_dqdPE4(Bit#(32) v);
    method Action a_curr_vec_in_AZ_dqdPE4(Bit#(32) v);
    method Action a_curr_vec_in_LX_dqdPE4(Bit#(32) v);
    method Action a_curr_vec_in_LY_dqdPE4(Bit#(32) v);
    method Action a_curr_vec_in_LZ_dqdPE4(Bit#(32) v);
    method Action a_curr_vec_in_AX_dqdPE5(Bit#(32) v);
    method Action a_curr_vec_in_AY_dqdPE5(Bit#(32) v);
    method Action a_curr_vec_in_AZ_dqdPE5(Bit#(32) v);
    method Action a_curr_vec_in_LX_dqdPE5(Bit#(32) v);
    method Action a_curr_vec_in_LY_dqdPE5(Bit#(32) v);
    method Action a_curr_vec_in_LZ_dqdPE5(Bit#(32) v);
    method Action a_curr_vec_in_AX_dqdPE6(Bit#(32) v);
    method Action a_curr_vec_in_AY_dqdPE6(Bit#(32) v);
    method Action a_curr_vec_in_AZ_dqdPE6(Bit#(32) v);
    method Action a_curr_vec_in_LX_dqdPE6(Bit#(32) v);
    method Action a_curr_vec_in_LY_dqdPE6(Bit#(32) v);
    method Action a_curr_vec_in_LZ_dqdPE6(Bit#(32) v);
    method Action a_curr_vec_in_AX_dqdPE7(Bit#(32) v);
    method Action a_curr_vec_in_AY_dqdPE7(Bit#(32) v);
    method Action a_curr_vec_in_AZ_dqdPE7(Bit#(32) v);
    method Action a_curr_vec_in_LX_dqdPE7(Bit#(32) v);
    method Action a_curr_vec_in_LY_dqdPE7(Bit#(32) v);
    method Action a_curr_vec_in_LZ_dqdPE7(Bit#(32) v);
    method Action v_prev_vec_in_AX_dqPE1(Bit#(32) v);
    method Action v_prev_vec_in_AY_dqPE1(Bit#(32) v);
    method Action v_prev_vec_in_AZ_dqPE1(Bit#(32) v);
    method Action v_prev_vec_in_LX_dqPE1(Bit#(32) v);
    method Action v_prev_vec_in_LY_dqPE1(Bit#(32) v);
    method Action v_prev_vec_in_LZ_dqPE1(Bit#(32) v);
    method Action v_prev_vec_in_AX_dqPE2(Bit#(32) v);
    method Action v_prev_vec_in_AY_dqPE2(Bit#(32) v);
    method Action v_prev_vec_in_AZ_dqPE2(Bit#(32) v);
    method Action v_prev_vec_in_LX_dqPE2(Bit#(32) v);
    method Action v_prev_vec_in_LY_dqPE2(Bit#(32) v);
    method Action v_prev_vec_in_LZ_dqPE2(Bit#(32) v);
    method Action v_prev_vec_in_AX_dqPE3(Bit#(32) v);
    method Action v_prev_vec_in_AY_dqPE3(Bit#(32) v);
    method Action v_prev_vec_in_AZ_dqPE3(Bit#(32) v);
    method Action v_prev_vec_in_LX_dqPE3(Bit#(32) v);
    method Action v_prev_vec_in_LY_dqPE3(Bit#(32) v);
    method Action v_prev_vec_in_LZ_dqPE3(Bit#(32) v);
    method Action v_prev_vec_in_AX_dqPE4(Bit#(32) v);
    method Action v_prev_vec_in_AY_dqPE4(Bit#(32) v);
    method Action v_prev_vec_in_AZ_dqPE4(Bit#(32) v);
    method Action v_prev_vec_in_LX_dqPE4(Bit#(32) v);
    method Action v_prev_vec_in_LY_dqPE4(Bit#(32) v);
    method Action v_prev_vec_in_LZ_dqPE4(Bit#(32) v);
    method Action v_prev_vec_in_AX_dqPE5(Bit#(32) v);
    method Action v_prev_vec_in_AY_dqPE5(Bit#(32) v);
    method Action v_prev_vec_in_AZ_dqPE5(Bit#(32) v);
    method Action v_prev_vec_in_LX_dqPE5(Bit#(32) v);
    method Action v_prev_vec_in_LY_dqPE5(Bit#(32) v);
    method Action v_prev_vec_in_LZ_dqPE5(Bit#(32) v);
    method Action v_prev_vec_in_AX_dqPE6(Bit#(32) v);
    method Action v_prev_vec_in_AY_dqPE6(Bit#(32) v);
    method Action v_prev_vec_in_AZ_dqPE6(Bit#(32) v);
    method Action v_prev_vec_in_LX_dqPE6(Bit#(32) v);
    method Action v_prev_vec_in_LY_dqPE6(Bit#(32) v);
    method Action v_prev_vec_in_LZ_dqPE6(Bit#(32) v);
    method Action v_prev_vec_in_AX_dqPE7(Bit#(32) v);
    method Action v_prev_vec_in_AY_dqPE7(Bit#(32) v);
    method Action v_prev_vec_in_AZ_dqPE7(Bit#(32) v);
    method Action v_prev_vec_in_LX_dqPE7(Bit#(32) v);
    method Action v_prev_vec_in_LY_dqPE7(Bit#(32) v);
    method Action v_prev_vec_in_LZ_dqPE7(Bit#(32) v);
    method Action a_prev_vec_in_AX_dqPE1(Bit#(32) v);
    method Action a_prev_vec_in_AY_dqPE1(Bit#(32) v);
    method Action a_prev_vec_in_AZ_dqPE1(Bit#(32) v);
    method Action a_prev_vec_in_LX_dqPE1(Bit#(32) v);
    method Action a_prev_vec_in_LY_dqPE1(Bit#(32) v);
    method Action a_prev_vec_in_LZ_dqPE1(Bit#(32) v);
    method Action a_prev_vec_in_AX_dqPE2(Bit#(32) v);
    method Action a_prev_vec_in_AY_dqPE2(Bit#(32) v);
    method Action a_prev_vec_in_AZ_dqPE2(Bit#(32) v);
    method Action a_prev_vec_in_LX_dqPE2(Bit#(32) v);
    method Action a_prev_vec_in_LY_dqPE2(Bit#(32) v);
    method Action a_prev_vec_in_LZ_dqPE2(Bit#(32) v);
    method Action a_prev_vec_in_AX_dqPE3(Bit#(32) v);
    method Action a_prev_vec_in_AY_dqPE3(Bit#(32) v);
    method Action a_prev_vec_in_AZ_dqPE3(Bit#(32) v);
    method Action a_prev_vec_in_LX_dqPE3(Bit#(32) v);
    method Action a_prev_vec_in_LY_dqPE3(Bit#(32) v);
    method Action a_prev_vec_in_LZ_dqPE3(Bit#(32) v);
    method Action a_prev_vec_in_AX_dqPE4(Bit#(32) v);
    method Action a_prev_vec_in_AY_dqPE4(Bit#(32) v);
    method Action a_prev_vec_in_AZ_dqPE4(Bit#(32) v);
    method Action a_prev_vec_in_LX_dqPE4(Bit#(32) v);
    method Action a_prev_vec_in_LY_dqPE4(Bit#(32) v);
    method Action a_prev_vec_in_LZ_dqPE4(Bit#(32) v);
    method Action a_prev_vec_in_AX_dqPE5(Bit#(32) v);
    method Action a_prev_vec_in_AY_dqPE5(Bit#(32) v);
    method Action a_prev_vec_in_AZ_dqPE5(Bit#(32) v);
    method Action a_prev_vec_in_LX_dqPE5(Bit#(32) v);
    method Action a_prev_vec_in_LY_dqPE5(Bit#(32) v);
    method Action a_prev_vec_in_LZ_dqPE5(Bit#(32) v);
    method Action a_prev_vec_in_AX_dqPE6(Bit#(32) v);
    method Action a_prev_vec_in_AY_dqPE6(Bit#(32) v);
    method Action a_prev_vec_in_AZ_dqPE6(Bit#(32) v);
    method Action a_prev_vec_in_LX_dqPE6(Bit#(32) v);
    method Action a_prev_vec_in_LY_dqPE6(Bit#(32) v);
    method Action a_prev_vec_in_LZ_dqPE6(Bit#(32) v);
    method Action a_prev_vec_in_AX_dqPE7(Bit#(32) v);
    method Action a_prev_vec_in_AY_dqPE7(Bit#(32) v);
    method Action a_prev_vec_in_AZ_dqPE7(Bit#(32) v);
    method Action a_prev_vec_in_LX_dqPE7(Bit#(32) v);
    method Action a_prev_vec_in_LY_dqPE7(Bit#(32) v);
    method Action a_prev_vec_in_LZ_dqPE7(Bit#(32) v);

    method Action dvdq_prev_vec_in_AX_dqPE1(Bit#(32) v);
    method Action dvdq_prev_vec_in_AY_dqPE1(Bit#(32) v);
    method Action dvdq_prev_vec_in_AZ_dqPE1(Bit#(32) v);
    method Action dvdq_prev_vec_in_LX_dqPE1(Bit#(32) v);
    method Action dvdq_prev_vec_in_LY_dqPE1(Bit#(32) v);
    method Action dvdq_prev_vec_in_LZ_dqPE1(Bit#(32) v);
    method Action dvdq_prev_vec_in_AX_dqPE2(Bit#(32) v);
    method Action dvdq_prev_vec_in_AY_dqPE2(Bit#(32) v);
    method Action dvdq_prev_vec_in_AZ_dqPE2(Bit#(32) v);
    method Action dvdq_prev_vec_in_LX_dqPE2(Bit#(32) v);
    method Action dvdq_prev_vec_in_LY_dqPE2(Bit#(32) v);
    method Action dvdq_prev_vec_in_LZ_dqPE2(Bit#(32) v);
    method Action dvdq_prev_vec_in_AX_dqPE3(Bit#(32) v);
    method Action dvdq_prev_vec_in_AY_dqPE3(Bit#(32) v);
    method Action dvdq_prev_vec_in_AZ_dqPE3(Bit#(32) v);
    method Action dvdq_prev_vec_in_LX_dqPE3(Bit#(32) v);
    method Action dvdq_prev_vec_in_LY_dqPE3(Bit#(32) v);
    method Action dvdq_prev_vec_in_LZ_dqPE3(Bit#(32) v);
    method Action dvdq_prev_vec_in_AX_dqPE4(Bit#(32) v);
    method Action dvdq_prev_vec_in_AY_dqPE4(Bit#(32) v);
    method Action dvdq_prev_vec_in_AZ_dqPE4(Bit#(32) v);
    method Action dvdq_prev_vec_in_LX_dqPE4(Bit#(32) v);
    method Action dvdq_prev_vec_in_LY_dqPE4(Bit#(32) v);
    method Action dvdq_prev_vec_in_LZ_dqPE4(Bit#(32) v);
    method Action dvdq_prev_vec_in_AX_dqPE5(Bit#(32) v);
    method Action dvdq_prev_vec_in_AY_dqPE5(Bit#(32) v);
    method Action dvdq_prev_vec_in_AZ_dqPE5(Bit#(32) v);
    method Action dvdq_prev_vec_in_LX_dqPE5(Bit#(32) v);
    method Action dvdq_prev_vec_in_LY_dqPE5(Bit#(32) v);
    method Action dvdq_prev_vec_in_LZ_dqPE5(Bit#(32) v);
    method Action dvdq_prev_vec_in_AX_dqPE6(Bit#(32) v);
    method Action dvdq_prev_vec_in_AY_dqPE6(Bit#(32) v);
    method Action dvdq_prev_vec_in_AZ_dqPE6(Bit#(32) v);
    method Action dvdq_prev_vec_in_LX_dqPE6(Bit#(32) v);
    method Action dvdq_prev_vec_in_LY_dqPE6(Bit#(32) v);
    method Action dvdq_prev_vec_in_LZ_dqPE6(Bit#(32) v);
    method Action dvdq_prev_vec_in_AX_dqPE7(Bit#(32) v);
    method Action dvdq_prev_vec_in_AY_dqPE7(Bit#(32) v);
    method Action dvdq_prev_vec_in_AZ_dqPE7(Bit#(32) v);
    method Action dvdq_prev_vec_in_LX_dqPE7(Bit#(32) v);
    method Action dvdq_prev_vec_in_LY_dqPE7(Bit#(32) v);
    method Action dvdq_prev_vec_in_LZ_dqPE7(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AX_dqdPE1(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AY_dqdPE1(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AZ_dqdPE1(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LX_dqdPE1(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LY_dqdPE1(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LZ_dqdPE1(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AX_dqdPE2(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AY_dqdPE2(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AZ_dqdPE2(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LX_dqdPE2(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LY_dqdPE2(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LZ_dqdPE2(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AX_dqdPE3(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AY_dqdPE3(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AZ_dqdPE3(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LX_dqdPE3(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LY_dqdPE3(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LZ_dqdPE3(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AX_dqdPE4(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AY_dqdPE4(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AZ_dqdPE4(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LX_dqdPE4(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LY_dqdPE4(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LZ_dqdPE4(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AX_dqdPE5(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AY_dqdPE5(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AZ_dqdPE5(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LX_dqdPE5(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LY_dqdPE5(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LZ_dqdPE5(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AX_dqdPE6(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AY_dqdPE6(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AZ_dqdPE6(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LX_dqdPE6(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LY_dqdPE6(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LZ_dqdPE6(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AX_dqdPE7(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AY_dqdPE7(Bit#(32) v);
    method Action dvdqd_prev_vec_in_AZ_dqdPE7(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LX_dqdPE7(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LY_dqdPE7(Bit#(32) v);
    method Action dvdqd_prev_vec_in_LZ_dqdPE7(Bit#(32) v);
    method Action dadq_prev_vec_in_AX_dqPE1(Bit#(32) v);
    method Action dadq_prev_vec_in_AY_dqPE1(Bit#(32) v);
    method Action dadq_prev_vec_in_AZ_dqPE1(Bit#(32) v);
    method Action dadq_prev_vec_in_LX_dqPE1(Bit#(32) v);
    method Action dadq_prev_vec_in_LY_dqPE1(Bit#(32) v);
    method Action dadq_prev_vec_in_LZ_dqPE1(Bit#(32) v);
    method Action dadq_prev_vec_in_AX_dqPE2(Bit#(32) v);
    method Action dadq_prev_vec_in_AY_dqPE2(Bit#(32) v);
    method Action dadq_prev_vec_in_AZ_dqPE2(Bit#(32) v);
    method Action dadq_prev_vec_in_LX_dqPE2(Bit#(32) v);
    method Action dadq_prev_vec_in_LY_dqPE2(Bit#(32) v);
    method Action dadq_prev_vec_in_LZ_dqPE2(Bit#(32) v);
    method Action dadq_prev_vec_in_AX_dqPE3(Bit#(32) v);
    method Action dadq_prev_vec_in_AY_dqPE3(Bit#(32) v);
    method Action dadq_prev_vec_in_AZ_dqPE3(Bit#(32) v);
    method Action dadq_prev_vec_in_LX_dqPE3(Bit#(32) v);
    method Action dadq_prev_vec_in_LY_dqPE3(Bit#(32) v);
    method Action dadq_prev_vec_in_LZ_dqPE3(Bit#(32) v);
    method Action dadq_prev_vec_in_AX_dqPE4(Bit#(32) v);
    method Action dadq_prev_vec_in_AY_dqPE4(Bit#(32) v);
    method Action dadq_prev_vec_in_AZ_dqPE4(Bit#(32) v);
    method Action dadq_prev_vec_in_LX_dqPE4(Bit#(32) v);
    method Action dadq_prev_vec_in_LY_dqPE4(Bit#(32) v);
    method Action dadq_prev_vec_in_LZ_dqPE4(Bit#(32) v);
    method Action dadq_prev_vec_in_AX_dqPE5(Bit#(32) v);
    method Action dadq_prev_vec_in_AY_dqPE5(Bit#(32) v);
    method Action dadq_prev_vec_in_AZ_dqPE5(Bit#(32) v);
    method Action dadq_prev_vec_in_LX_dqPE5(Bit#(32) v);
    method Action dadq_prev_vec_in_LY_dqPE5(Bit#(32) v);
    method Action dadq_prev_vec_in_LZ_dqPE5(Bit#(32) v);
    method Action dadq_prev_vec_in_AX_dqPE6(Bit#(32) v);
    method Action dadq_prev_vec_in_AY_dqPE6(Bit#(32) v);
    method Action dadq_prev_vec_in_AZ_dqPE6(Bit#(32) v);
    method Action dadq_prev_vec_in_LX_dqPE6(Bit#(32) v);
    method Action dadq_prev_vec_in_LY_dqPE6(Bit#(32) v);
    method Action dadq_prev_vec_in_LZ_dqPE6(Bit#(32) v);
    method Action dadq_prev_vec_in_AX_dqPE7(Bit#(32) v);
    method Action dadq_prev_vec_in_AY_dqPE7(Bit#(32) v);
    method Action dadq_prev_vec_in_AZ_dqPE7(Bit#(32) v);
    method Action dadq_prev_vec_in_LX_dqPE7(Bit#(32) v);
    method Action dadq_prev_vec_in_LY_dqPE7(Bit#(32) v);
    method Action dadq_prev_vec_in_LZ_dqPE7(Bit#(32) v);
    method Action dadqd_prev_vec_in_AX_dqdPE1(Bit#(32) v);
    method Action dadqd_prev_vec_in_AY_dqdPE1(Bit#(32) v);
    method Action dadqd_prev_vec_in_AZ_dqdPE1(Bit#(32) v);
    method Action dadqd_prev_vec_in_LX_dqdPE1(Bit#(32) v);
    method Action dadqd_prev_vec_in_LY_dqdPE1(Bit#(32) v);
    method Action dadqd_prev_vec_in_LZ_dqdPE1(Bit#(32) v);
    method Action dadqd_prev_vec_in_AX_dqdPE2(Bit#(32) v);
    method Action dadqd_prev_vec_in_AY_dqdPE2(Bit#(32) v);
    method Action dadqd_prev_vec_in_AZ_dqdPE2(Bit#(32) v);
    method Action dadqd_prev_vec_in_LX_dqdPE2(Bit#(32) v);
    method Action dadqd_prev_vec_in_LY_dqdPE2(Bit#(32) v);
    method Action dadqd_prev_vec_in_LZ_dqdPE2(Bit#(32) v);
    method Action dadqd_prev_vec_in_AX_dqdPE3(Bit#(32) v);
    method Action dadqd_prev_vec_in_AY_dqdPE3(Bit#(32) v);
    method Action dadqd_prev_vec_in_AZ_dqdPE3(Bit#(32) v);
    method Action dadqd_prev_vec_in_LX_dqdPE3(Bit#(32) v);
    method Action dadqd_prev_vec_in_LY_dqdPE3(Bit#(32) v);
    method Action dadqd_prev_vec_in_LZ_dqdPE3(Bit#(32) v);
    method Action dadqd_prev_vec_in_AX_dqdPE4(Bit#(32) v);
    method Action dadqd_prev_vec_in_AY_dqdPE4(Bit#(32) v);
    method Action dadqd_prev_vec_in_AZ_dqdPE4(Bit#(32) v);
    method Action dadqd_prev_vec_in_LX_dqdPE4(Bit#(32) v);
    method Action dadqd_prev_vec_in_LY_dqdPE4(Bit#(32) v);
    method Action dadqd_prev_vec_in_LZ_dqdPE4(Bit#(32) v);
    method Action dadqd_prev_vec_in_AX_dqdPE5(Bit#(32) v);
    method Action dadqd_prev_vec_in_AY_dqdPE5(Bit#(32) v);
    method Action dadqd_prev_vec_in_AZ_dqdPE5(Bit#(32) v);
    method Action dadqd_prev_vec_in_LX_dqdPE5(Bit#(32) v);
    method Action dadqd_prev_vec_in_LY_dqdPE5(Bit#(32) v);
    method Action dadqd_prev_vec_in_LZ_dqdPE5(Bit#(32) v);
    method Action dadqd_prev_vec_in_AX_dqdPE6(Bit#(32) v);
    method Action dadqd_prev_vec_in_AY_dqdPE6(Bit#(32) v);
    method Action dadqd_prev_vec_in_AZ_dqdPE6(Bit#(32) v);
    method Action dadqd_prev_vec_in_LX_dqdPE6(Bit#(32) v);
    method Action dadqd_prev_vec_in_LY_dqdPE6(Bit#(32) v);
    method Action dadqd_prev_vec_in_LZ_dqdPE6(Bit#(32) v);
    method Action dadqd_prev_vec_in_AX_dqdPE7(Bit#(32) v);
    method Action dadqd_prev_vec_in_AY_dqdPE7(Bit#(32) v);
    method Action dadqd_prev_vec_in_AZ_dqdPE7(Bit#(32) v);
    method Action dadqd_prev_vec_in_LX_dqdPE7(Bit#(32) v);
    method Action dadqd_prev_vec_in_LY_dqdPE7(Bit#(32) v);
    method Action dadqd_prev_vec_in_LZ_dqdPE7(Bit#(32) v);

    //--------------------------

    // output_ready
    method Bit#(1) output_ready();

    //-------- RNEA OUTPUTS -----

    method Bit#(32) v_curr_vec_out_AX_rnea();
    method Bit#(32) v_curr_vec_out_AY_rnea();
    method Bit#(32) v_curr_vec_out_AZ_rnea();
    method Bit#(32) v_curr_vec_out_LX_rnea();
    method Bit#(32) v_curr_vec_out_LY_rnea();
    method Bit#(32) v_curr_vec_out_LZ_rnea();
    method Bit#(32) a_curr_vec_out_AX_rnea();
    method Bit#(32) a_curr_vec_out_AY_rnea();
    method Bit#(32) a_curr_vec_out_AZ_rnea();
    method Bit#(32) a_curr_vec_out_LX_rnea();
    method Bit#(32) a_curr_vec_out_LY_rnea();
    method Bit#(32) a_curr_vec_out_LZ_rnea();
    method Bit#(32) f_curr_vec_out_AX_rnea();
    method Bit#(32) f_curr_vec_out_AY_rnea();
    method Bit#(32) f_curr_vec_out_AZ_rnea();
    method Bit#(32) f_curr_vec_out_LX_rnea();
    method Bit#(32) f_curr_vec_out_LY_rnea();
    method Bit#(32) f_curr_vec_out_LZ_rnea();

    //-----------------------

    //----------- DQ DQD OUTPUTS -----

    method Bit#(32) dfdq_curr_vec_out_AX_dqPE1();
    method Bit#(32) dfdq_curr_vec_out_AY_dqPE1();
    method Bit#(32) dfdq_curr_vec_out_AZ_dqPE1();
    method Bit#(32) dfdq_curr_vec_out_LX_dqPE1();
    method Bit#(32) dfdq_curr_vec_out_LY_dqPE1();
    method Bit#(32) dfdq_curr_vec_out_LZ_dqPE1();
    method Bit#(32) dfdq_curr_vec_out_AX_dqPE2();
    method Bit#(32) dfdq_curr_vec_out_AY_dqPE2();
    method Bit#(32) dfdq_curr_vec_out_AZ_dqPE2();
    method Bit#(32) dfdq_curr_vec_out_LX_dqPE2();
    method Bit#(32) dfdq_curr_vec_out_LY_dqPE2();
    method Bit#(32) dfdq_curr_vec_out_LZ_dqPE2();
    method Bit#(32) dfdq_curr_vec_out_AX_dqPE3();
    method Bit#(32) dfdq_curr_vec_out_AY_dqPE3();
    method Bit#(32) dfdq_curr_vec_out_AZ_dqPE3();
    method Bit#(32) dfdq_curr_vec_out_LX_dqPE3();
    method Bit#(32) dfdq_curr_vec_out_LY_dqPE3();
    method Bit#(32) dfdq_curr_vec_out_LZ_dqPE3();
    method Bit#(32) dfdq_curr_vec_out_AX_dqPE4();
    method Bit#(32) dfdq_curr_vec_out_AY_dqPE4();
    method Bit#(32) dfdq_curr_vec_out_AZ_dqPE4();
    method Bit#(32) dfdq_curr_vec_out_LX_dqPE4();
    method Bit#(32) dfdq_curr_vec_out_LY_dqPE4();
    method Bit#(32) dfdq_curr_vec_out_LZ_dqPE4();
    method Bit#(32) dfdq_curr_vec_out_AX_dqPE5();
    method Bit#(32) dfdq_curr_vec_out_AY_dqPE5();
    method Bit#(32) dfdq_curr_vec_out_AZ_dqPE5();
    method Bit#(32) dfdq_curr_vec_out_LX_dqPE5();
    method Bit#(32) dfdq_curr_vec_out_LY_dqPE5();
    method Bit#(32) dfdq_curr_vec_out_LZ_dqPE5();
    method Bit#(32) dfdq_curr_vec_out_AX_dqPE6();
    method Bit#(32) dfdq_curr_vec_out_AY_dqPE6();
    method Bit#(32) dfdq_curr_vec_out_AZ_dqPE6();
    method Bit#(32) dfdq_curr_vec_out_LX_dqPE6();
    method Bit#(32) dfdq_curr_vec_out_LY_dqPE6();
    method Bit#(32) dfdq_curr_vec_out_LZ_dqPE6();
    method Bit#(32) dfdq_curr_vec_out_AX_dqPE7();
    method Bit#(32) dfdq_curr_vec_out_AY_dqPE7();
    method Bit#(32) dfdq_curr_vec_out_AZ_dqPE7();
    method Bit#(32) dfdq_curr_vec_out_LX_dqPE7();
    method Bit#(32) dfdq_curr_vec_out_LY_dqPE7();
    method Bit#(32) dfdq_curr_vec_out_LZ_dqPE7();
    method Bit#(32) dfdqd_curr_vec_out_AX_dqdPE1();
    method Bit#(32) dfdqd_curr_vec_out_AY_dqdPE1();
    method Bit#(32) dfdqd_curr_vec_out_AZ_dqdPE1();
    method Bit#(32) dfdqd_curr_vec_out_LX_dqdPE1();
    method Bit#(32) dfdqd_curr_vec_out_LY_dqdPE1();
    method Bit#(32) dfdqd_curr_vec_out_LZ_dqdPE1();
    method Bit#(32) dfdqd_curr_vec_out_AX_dqdPE2();
    method Bit#(32) dfdqd_curr_vec_out_AY_dqdPE2();
    method Bit#(32) dfdqd_curr_vec_out_AZ_dqdPE2();
    method Bit#(32) dfdqd_curr_vec_out_LX_dqdPE2();
    method Bit#(32) dfdqd_curr_vec_out_LY_dqdPE2();
    method Bit#(32) dfdqd_curr_vec_out_LZ_dqdPE2();
    method Bit#(32) dfdqd_curr_vec_out_AX_dqdPE3();
    method Bit#(32) dfdqd_curr_vec_out_AY_dqdPE3();
    method Bit#(32) dfdqd_curr_vec_out_AZ_dqdPE3();
    method Bit#(32) dfdqd_curr_vec_out_LX_dqdPE3();
    method Bit#(32) dfdqd_curr_vec_out_LY_dqdPE3();
    method Bit#(32) dfdqd_curr_vec_out_LZ_dqdPE3();
    method Bit#(32) dfdqd_curr_vec_out_AX_dqdPE4();
    method Bit#(32) dfdqd_curr_vec_out_AY_dqdPE4();
    method Bit#(32) dfdqd_curr_vec_out_AZ_dqdPE4();
    method Bit#(32) dfdqd_curr_vec_out_LX_dqdPE4();
    method Bit#(32) dfdqd_curr_vec_out_LY_dqdPE4();
    method Bit#(32) dfdqd_curr_vec_out_LZ_dqdPE4();
    method Bit#(32) dfdqd_curr_vec_out_AX_dqdPE5();
    method Bit#(32) dfdqd_curr_vec_out_AY_dqdPE5();
    method Bit#(32) dfdqd_curr_vec_out_AZ_dqdPE5();
    method Bit#(32) dfdqd_curr_vec_out_LX_dqdPE5();
    method Bit#(32) dfdqd_curr_vec_out_LY_dqdPE5();
    method Bit#(32) dfdqd_curr_vec_out_LZ_dqdPE5();
    method Bit#(32) dfdqd_curr_vec_out_AX_dqdPE6();
    method Bit#(32) dfdqd_curr_vec_out_AY_dqdPE6();
    method Bit#(32) dfdqd_curr_vec_out_AZ_dqdPE6();
    method Bit#(32) dfdqd_curr_vec_out_LX_dqdPE6();
    method Bit#(32) dfdqd_curr_vec_out_LY_dqdPE6();
    method Bit#(32) dfdqd_curr_vec_out_LZ_dqdPE6();
    method Bit#(32) dfdqd_curr_vec_out_AX_dqdPE7();
    method Bit#(32) dfdqd_curr_vec_out_AY_dqdPE7();
    method Bit#(32) dfdqd_curr_vec_out_AZ_dqdPE7();
    method Bit#(32) dfdqd_curr_vec_out_LX_dqdPE7();
    method Bit#(32) dfdqd_curr_vec_out_LY_dqdPE7();
    method Bit#(32) dfdqd_curr_vec_out_LZ_dqdPE7();

    method Bit#(32) dvdq_curr_vec_out_AX_dqPE1();
    method Bit#(32) dvdq_curr_vec_out_AY_dqPE1();
    method Bit#(32) dvdq_curr_vec_out_AZ_dqPE1();
    method Bit#(32) dvdq_curr_vec_out_LX_dqPE1();
    method Bit#(32) dvdq_curr_vec_out_LY_dqPE1();
    method Bit#(32) dvdq_curr_vec_out_LZ_dqPE1();
    method Bit#(32) dvdq_curr_vec_out_AX_dqPE2();
    method Bit#(32) dvdq_curr_vec_out_AY_dqPE2();
    method Bit#(32) dvdq_curr_vec_out_AZ_dqPE2();
    method Bit#(32) dvdq_curr_vec_out_LX_dqPE2();
    method Bit#(32) dvdq_curr_vec_out_LY_dqPE2();
    method Bit#(32) dvdq_curr_vec_out_LZ_dqPE2();
    method Bit#(32) dvdq_curr_vec_out_AX_dqPE3();
    method Bit#(32) dvdq_curr_vec_out_AY_dqPE3();
    method Bit#(32) dvdq_curr_vec_out_AZ_dqPE3();
    method Bit#(32) dvdq_curr_vec_out_LX_dqPE3();
    method Bit#(32) dvdq_curr_vec_out_LY_dqPE3();
    method Bit#(32) dvdq_curr_vec_out_LZ_dqPE3();
    method Bit#(32) dvdq_curr_vec_out_AX_dqPE4();
    method Bit#(32) dvdq_curr_vec_out_AY_dqPE4();
    method Bit#(32) dvdq_curr_vec_out_AZ_dqPE4();
    method Bit#(32) dvdq_curr_vec_out_LX_dqPE4();
    method Bit#(32) dvdq_curr_vec_out_LY_dqPE4();
    method Bit#(32) dvdq_curr_vec_out_LZ_dqPE4();
    method Bit#(32) dvdq_curr_vec_out_AX_dqPE5();
    method Bit#(32) dvdq_curr_vec_out_AY_dqPE5();
    method Bit#(32) dvdq_curr_vec_out_AZ_dqPE5();
    method Bit#(32) dvdq_curr_vec_out_LX_dqPE5();
    method Bit#(32) dvdq_curr_vec_out_LY_dqPE5();
    method Bit#(32) dvdq_curr_vec_out_LZ_dqPE5();
    method Bit#(32) dvdq_curr_vec_out_AX_dqPE6();
    method Bit#(32) dvdq_curr_vec_out_AY_dqPE6();
    method Bit#(32) dvdq_curr_vec_out_AZ_dqPE6();
    method Bit#(32) dvdq_curr_vec_out_LX_dqPE6();
    method Bit#(32) dvdq_curr_vec_out_LY_dqPE6();
    method Bit#(32) dvdq_curr_vec_out_LZ_dqPE6();
    method Bit#(32) dvdq_curr_vec_out_AX_dqPE7();
    method Bit#(32) dvdq_curr_vec_out_AY_dqPE7();
    method Bit#(32) dvdq_curr_vec_out_AZ_dqPE7();
    method Bit#(32) dvdq_curr_vec_out_LX_dqPE7();
    method Bit#(32) dvdq_curr_vec_out_LY_dqPE7();
    method Bit#(32) dvdq_curr_vec_out_LZ_dqPE7();
    method Bit#(32) dvdqd_curr_vec_out_AX_dqdPE1();
    method Bit#(32) dvdqd_curr_vec_out_AY_dqdPE1();
    method Bit#(32) dvdqd_curr_vec_out_AZ_dqdPE1();
    method Bit#(32) dvdqd_curr_vec_out_LX_dqdPE1();
    method Bit#(32) dvdqd_curr_vec_out_LY_dqdPE1();
    method Bit#(32) dvdqd_curr_vec_out_LZ_dqdPE1();
    method Bit#(32) dvdqd_curr_vec_out_AX_dqdPE2();
    method Bit#(32) dvdqd_curr_vec_out_AY_dqdPE2();
    method Bit#(32) dvdqd_curr_vec_out_AZ_dqdPE2();
    method Bit#(32) dvdqd_curr_vec_out_LX_dqdPE2();
    method Bit#(32) dvdqd_curr_vec_out_LY_dqdPE2();
    method Bit#(32) dvdqd_curr_vec_out_LZ_dqdPE2();
    method Bit#(32) dvdqd_curr_vec_out_AX_dqdPE3();
    method Bit#(32) dvdqd_curr_vec_out_AY_dqdPE3();
    method Bit#(32) dvdqd_curr_vec_out_AZ_dqdPE3();
    method Bit#(32) dvdqd_curr_vec_out_LX_dqdPE3();
    method Bit#(32) dvdqd_curr_vec_out_LY_dqdPE3();
    method Bit#(32) dvdqd_curr_vec_out_LZ_dqdPE3();
    method Bit#(32) dvdqd_curr_vec_out_AX_dqdPE4();
    method Bit#(32) dvdqd_curr_vec_out_AY_dqdPE4();
    method Bit#(32) dvdqd_curr_vec_out_AZ_dqdPE4();
    method Bit#(32) dvdqd_curr_vec_out_LX_dqdPE4();
    method Bit#(32) dvdqd_curr_vec_out_LY_dqdPE4();
    method Bit#(32) dvdqd_curr_vec_out_LZ_dqdPE4();
    method Bit#(32) dvdqd_curr_vec_out_AX_dqdPE5();
    method Bit#(32) dvdqd_curr_vec_out_AY_dqdPE5();
    method Bit#(32) dvdqd_curr_vec_out_AZ_dqdPE5();
    method Bit#(32) dvdqd_curr_vec_out_LX_dqdPE5();
    method Bit#(32) dvdqd_curr_vec_out_LY_dqdPE5();
    method Bit#(32) dvdqd_curr_vec_out_LZ_dqdPE5();
    method Bit#(32) dvdqd_curr_vec_out_AX_dqdPE6();
    method Bit#(32) dvdqd_curr_vec_out_AY_dqdPE6();
    method Bit#(32) dvdqd_curr_vec_out_AZ_dqdPE6();
    method Bit#(32) dvdqd_curr_vec_out_LX_dqdPE6();
    method Bit#(32) dvdqd_curr_vec_out_LY_dqdPE6();
    method Bit#(32) dvdqd_curr_vec_out_LZ_dqdPE6();
    method Bit#(32) dvdqd_curr_vec_out_AX_dqdPE7();
    method Bit#(32) dvdqd_curr_vec_out_AY_dqdPE7();
    method Bit#(32) dvdqd_curr_vec_out_AZ_dqdPE7();
    method Bit#(32) dvdqd_curr_vec_out_LX_dqdPE7();
    method Bit#(32) dvdqd_curr_vec_out_LY_dqdPE7();
    method Bit#(32) dvdqd_curr_vec_out_LZ_dqdPE7();
    method Bit#(32) dadq_curr_vec_out_AX_dqPE1();
    method Bit#(32) dadq_curr_vec_out_AY_dqPE1();
    method Bit#(32) dadq_curr_vec_out_AZ_dqPE1();
    method Bit#(32) dadq_curr_vec_out_LX_dqPE1();
    method Bit#(32) dadq_curr_vec_out_LY_dqPE1();
    method Bit#(32) dadq_curr_vec_out_LZ_dqPE1();
    method Bit#(32) dadq_curr_vec_out_AX_dqPE2();
    method Bit#(32) dadq_curr_vec_out_AY_dqPE2();
    method Bit#(32) dadq_curr_vec_out_AZ_dqPE2();
    method Bit#(32) dadq_curr_vec_out_LX_dqPE2();
    method Bit#(32) dadq_curr_vec_out_LY_dqPE2();
    method Bit#(32) dadq_curr_vec_out_LZ_dqPE2();
    method Bit#(32) dadq_curr_vec_out_AX_dqPE3();
    method Bit#(32) dadq_curr_vec_out_AY_dqPE3();
    method Bit#(32) dadq_curr_vec_out_AZ_dqPE3();
    method Bit#(32) dadq_curr_vec_out_LX_dqPE3();
    method Bit#(32) dadq_curr_vec_out_LY_dqPE3();
    method Bit#(32) dadq_curr_vec_out_LZ_dqPE3();
    method Bit#(32) dadq_curr_vec_out_AX_dqPE4();
    method Bit#(32) dadq_curr_vec_out_AY_dqPE4();
    method Bit#(32) dadq_curr_vec_out_AZ_dqPE4();
    method Bit#(32) dadq_curr_vec_out_LX_dqPE4();
    method Bit#(32) dadq_curr_vec_out_LY_dqPE4();
    method Bit#(32) dadq_curr_vec_out_LZ_dqPE4();
    method Bit#(32) dadq_curr_vec_out_AX_dqPE5();
    method Bit#(32) dadq_curr_vec_out_AY_dqPE5();
    method Bit#(32) dadq_curr_vec_out_AZ_dqPE5();
    method Bit#(32) dadq_curr_vec_out_LX_dqPE5();
    method Bit#(32) dadq_curr_vec_out_LY_dqPE5();
    method Bit#(32) dadq_curr_vec_out_LZ_dqPE5();
    method Bit#(32) dadq_curr_vec_out_AX_dqPE6();
    method Bit#(32) dadq_curr_vec_out_AY_dqPE6();
    method Bit#(32) dadq_curr_vec_out_AZ_dqPE6();
    method Bit#(32) dadq_curr_vec_out_LX_dqPE6();
    method Bit#(32) dadq_curr_vec_out_LY_dqPE6();
    method Bit#(32) dadq_curr_vec_out_LZ_dqPE6();
    method Bit#(32) dadq_curr_vec_out_AX_dqPE7();
    method Bit#(32) dadq_curr_vec_out_AY_dqPE7();
    method Bit#(32) dadq_curr_vec_out_AZ_dqPE7();
    method Bit#(32) dadq_curr_vec_out_LX_dqPE7();
    method Bit#(32) dadq_curr_vec_out_LY_dqPE7();
    method Bit#(32) dadq_curr_vec_out_LZ_dqPE7();
    method Bit#(32) dadqd_curr_vec_out_AX_dqdPE1();
    method Bit#(32) dadqd_curr_vec_out_AY_dqdPE1();
    method Bit#(32) dadqd_curr_vec_out_AZ_dqdPE1();
    method Bit#(32) dadqd_curr_vec_out_LX_dqdPE1();
    method Bit#(32) dadqd_curr_vec_out_LY_dqdPE1();
    method Bit#(32) dadqd_curr_vec_out_LZ_dqdPE1();
    method Bit#(32) dadqd_curr_vec_out_AX_dqdPE2();
    method Bit#(32) dadqd_curr_vec_out_AY_dqdPE2();
    method Bit#(32) dadqd_curr_vec_out_AZ_dqdPE2();
    method Bit#(32) dadqd_curr_vec_out_LX_dqdPE2();
    method Bit#(32) dadqd_curr_vec_out_LY_dqdPE2();
    method Bit#(32) dadqd_curr_vec_out_LZ_dqdPE2();
    method Bit#(32) dadqd_curr_vec_out_AX_dqdPE3();
    method Bit#(32) dadqd_curr_vec_out_AY_dqdPE3();
    method Bit#(32) dadqd_curr_vec_out_AZ_dqdPE3();
    method Bit#(32) dadqd_curr_vec_out_LX_dqdPE3();
    method Bit#(32) dadqd_curr_vec_out_LY_dqdPE3();
    method Bit#(32) dadqd_curr_vec_out_LZ_dqdPE3();
    method Bit#(32) dadqd_curr_vec_out_AX_dqdPE4();
    method Bit#(32) dadqd_curr_vec_out_AY_dqdPE4();
    method Bit#(32) dadqd_curr_vec_out_AZ_dqdPE4();
    method Bit#(32) dadqd_curr_vec_out_LX_dqdPE4();
    method Bit#(32) dadqd_curr_vec_out_LY_dqdPE4();
    method Bit#(32) dadqd_curr_vec_out_LZ_dqdPE4();
    method Bit#(32) dadqd_curr_vec_out_AX_dqdPE5();
    method Bit#(32) dadqd_curr_vec_out_AY_dqdPE5();
    method Bit#(32) dadqd_curr_vec_out_AZ_dqdPE5();
    method Bit#(32) dadqd_curr_vec_out_LX_dqdPE5();
    method Bit#(32) dadqd_curr_vec_out_LY_dqdPE5();
    method Bit#(32) dadqd_curr_vec_out_LZ_dqdPE5();
    method Bit#(32) dadqd_curr_vec_out_AX_dqdPE6();
    method Bit#(32) dadqd_curr_vec_out_AY_dqdPE6();
    method Bit#(32) dadqd_curr_vec_out_AZ_dqdPE6();
    method Bit#(32) dadqd_curr_vec_out_LX_dqdPE6();
    method Bit#(32) dadqd_curr_vec_out_LY_dqdPE6();
    method Bit#(32) dadqd_curr_vec_out_LZ_dqdPE6();
    method Bit#(32) dadqd_curr_vec_out_AX_dqdPE7();
    method Bit#(32) dadqd_curr_vec_out_AY_dqdPE7();
    method Bit#(32) dadqd_curr_vec_out_AZ_dqdPE7();
    method Bit#(32) dadqd_curr_vec_out_LX_dqdPE7();
    method Bit#(32) dadqd_curr_vec_out_LY_dqdPE7();
    method Bit#(32) dadqd_curr_vec_out_LZ_dqdPE7();

    //-----------------------

endinterface

import "BVI" fproc =
module mkFProc(FProc);
    default_clock clk();
    default_reset rst();
    input_clock (clk) <- exposeCurrentClock; 
    input_reset (reset) <- invertCurrentReset;
    method get_data() enable(get_data);

    method link_in_rnea(link_in_rnea) enable((*inhigh*) EN_link_in_rnea) ;
    method sinq_val_in_rnea(sinq_val_in_rnea) enable((*inhigh*) EN_sinq_val_in_rnea) ;
    method cosq_val_in_rnea(cosq_val_in_rnea) enable((*inhigh*) EN_cosq_val_in_rnea) ;
    method qd_val_in_rnea(qd_val_in_rnea) enable((*inhigh*) EN_qd_val_in_rnea) ;
    method qdd_val_in_rnea(qdd_val_in_rnea) enable((*inhigh*) EN_qdd_val_in_rnea) ;

    method v_prev_vec_in_AX_rnea(v_prev_vec_in_AX_rnea) enable((*inhigh*) EN_v_prev_vec_in_AX_rnea) ;
    method v_prev_vec_in_AY_rnea(v_prev_vec_in_AY_rnea) enable((*inhigh*) EN_v_prev_vec_in_AY_rnea) ;
    method v_prev_vec_in_AZ_rnea(v_prev_vec_in_AZ_rnea) enable((*inhigh*) EN_v_prev_vec_in_AZ_rnea) ;
    method v_prev_vec_in_LX_rnea(v_prev_vec_in_LX_rnea) enable((*inhigh*) EN_v_prev_vec_in_LX_rnea) ;
    method v_prev_vec_in_LY_rnea(v_prev_vec_in_LY_rnea) enable((*inhigh*) EN_v_prev_vec_in_LY_rnea) ;
    method v_prev_vec_in_LZ_rnea(v_prev_vec_in_LZ_rnea) enable((*inhigh*) EN_v_prev_vec_in_LZ_rnea) ;
    method a_prev_vec_in_AX_rnea(a_prev_vec_in_AX_rnea) enable((*inhigh*) EN_a_prev_vec_in_AX_rnea) ;
    method a_prev_vec_in_AY_rnea(a_prev_vec_in_AY_rnea) enable((*inhigh*) EN_a_prev_vec_in_AY_rnea) ;
    method a_prev_vec_in_AZ_rnea(a_prev_vec_in_AZ_rnea) enable((*inhigh*) EN_a_prev_vec_in_AZ_rnea) ;
    method a_prev_vec_in_LX_rnea(a_prev_vec_in_LX_rnea) enable((*inhigh*) EN_a_prev_vec_in_LX_rnea) ;
    method a_prev_vec_in_LY_rnea(a_prev_vec_in_LY_rnea) enable((*inhigh*) EN_a_prev_vec_in_LY_rnea) ;
    method a_prev_vec_in_LZ_rnea(a_prev_vec_in_LZ_rnea) enable((*inhigh*) EN_a_prev_vec_in_LZ_rnea) ;

    method link_in_dqPE1(link_in_dqPE1) enable((*inhigh*) EN_link_in_dqPE1) ;
    method link_in_dqPE2(link_in_dqPE2) enable((*inhigh*) EN_link_in_dqPE2) ;
    method link_in_dqPE3(link_in_dqPE3) enable((*inhigh*) EN_link_in_dqPE3) ;
    method link_in_dqPE4(link_in_dqPE4) enable((*inhigh*) EN_link_in_dqPE4) ;
    method link_in_dqPE5(link_in_dqPE5) enable((*inhigh*) EN_link_in_dqPE5) ;
    method link_in_dqPE6(link_in_dqPE6) enable((*inhigh*) EN_link_in_dqPE6) ;
    method link_in_dqPE7(link_in_dqPE7) enable((*inhigh*) EN_link_in_dqPE7) ;
    method link_in_dqdPE1(link_in_dqdPE1) enable((*inhigh*) EN_link_in_dqdPE1) ;
    method link_in_dqdPE2(link_in_dqdPE2) enable((*inhigh*) EN_link_in_dqdPE2) ;
    method link_in_dqdPE3(link_in_dqdPE3) enable((*inhigh*) EN_link_in_dqdPE3) ;
    method link_in_dqdPE4(link_in_dqdPE4) enable((*inhigh*) EN_link_in_dqdPE4) ;
    method link_in_dqdPE5(link_in_dqdPE5) enable((*inhigh*) EN_link_in_dqdPE5) ;
    method link_in_dqdPE6(link_in_dqdPE6) enable((*inhigh*) EN_link_in_dqdPE6) ;
    method link_in_dqdPE7(link_in_dqdPE7) enable((*inhigh*) EN_link_in_dqdPE7) ;
    method derv_in_dqPE1(derv_in_dqPE1) enable((*inhigh*) EN_derv_in_dqPE1) ;
    method derv_in_dqPE2(derv_in_dqPE2) enable((*inhigh*) EN_derv_in_dqPE2) ;
    method derv_in_dqPE3(derv_in_dqPE3) enable((*inhigh*) EN_derv_in_dqPE3) ;
    method derv_in_dqPE4(derv_in_dqPE4) enable((*inhigh*) EN_derv_in_dqPE4) ;
    method derv_in_dqPE5(derv_in_dqPE5) enable((*inhigh*) EN_derv_in_dqPE5) ;
    method derv_in_dqPE6(derv_in_dqPE6) enable((*inhigh*) EN_derv_in_dqPE6) ;
    method derv_in_dqPE7(derv_in_dqPE7) enable((*inhigh*) EN_derv_in_dqPE7) ;
    method derv_in_dqdPE1(derv_in_dqdPE1) enable((*inhigh*) EN_derv_in_dqdPE1) ;
    method derv_in_dqdPE2(derv_in_dqdPE2) enable((*inhigh*) EN_derv_in_dqdPE2) ;
    method derv_in_dqdPE3(derv_in_dqdPE3) enable((*inhigh*) EN_derv_in_dqdPE3) ;
    method derv_in_dqdPE4(derv_in_dqdPE4) enable((*inhigh*) EN_derv_in_dqdPE4) ;
    method derv_in_dqdPE5(derv_in_dqdPE5) enable((*inhigh*) EN_derv_in_dqdPE5) ;
    method derv_in_dqdPE6(derv_in_dqdPE6) enable((*inhigh*) EN_derv_in_dqdPE6) ;
    method derv_in_dqdPE7(derv_in_dqdPE7) enable((*inhigh*) EN_derv_in_dqdPE7) ;

    method sinq_val_in_dqPE1(sinq_val_in_dqPE1) enable((*inhigh*) EN_sinq_val_in_dqPE1) ;
    method sinq_val_in_dqPE2(sinq_val_in_dqPE2) enable((*inhigh*) EN_sinq_val_in_dqPE2) ;
    method sinq_val_in_dqPE3(sinq_val_in_dqPE3) enable((*inhigh*) EN_sinq_val_in_dqPE3) ;
    method sinq_val_in_dqPE4(sinq_val_in_dqPE4) enable((*inhigh*) EN_sinq_val_in_dqPE4) ;
    method sinq_val_in_dqPE5(sinq_val_in_dqPE5) enable((*inhigh*) EN_sinq_val_in_dqPE5) ;
    method sinq_val_in_dqPE6(sinq_val_in_dqPE6) enable((*inhigh*) EN_sinq_val_in_dqPE6) ;
    method sinq_val_in_dqPE7(sinq_val_in_dqPE7) enable((*inhigh*) EN_sinq_val_in_dqPE7) ;
    method sinq_val_in_dqdPE1(sinq_val_in_dqdPE1) enable((*inhigh*) EN_sinq_val_in_dqdPE1) ;
    method sinq_val_in_dqdPE2(sinq_val_in_dqdPE2) enable((*inhigh*) EN_sinq_val_in_dqdPE2) ;
    method sinq_val_in_dqdPE3(sinq_val_in_dqdPE3) enable((*inhigh*) EN_sinq_val_in_dqdPE3) ;
    method sinq_val_in_dqdPE4(sinq_val_in_dqdPE4) enable((*inhigh*) EN_sinq_val_in_dqdPE4) ;
    method sinq_val_in_dqdPE5(sinq_val_in_dqdPE5) enable((*inhigh*) EN_sinq_val_in_dqdPE5) ;
    method sinq_val_in_dqdPE6(sinq_val_in_dqdPE6) enable((*inhigh*) EN_sinq_val_in_dqdPE6) ;
    method sinq_val_in_dqdPE7(sinq_val_in_dqdPE7) enable((*inhigh*) EN_sinq_val_in_dqdPE7) ;
    method cosq_val_in_dqPE1(cosq_val_in_dqPE1) enable((*inhigh*) EN_cosq_val_in_dqPE1) ;
    method cosq_val_in_dqPE2(cosq_val_in_dqPE2) enable((*inhigh*) EN_cosq_val_in_dqPE2) ;
    method cosq_val_in_dqPE3(cosq_val_in_dqPE3) enable((*inhigh*) EN_cosq_val_in_dqPE3) ;
    method cosq_val_in_dqPE4(cosq_val_in_dqPE4) enable((*inhigh*) EN_cosq_val_in_dqPE4) ;
    method cosq_val_in_dqPE5(cosq_val_in_dqPE5) enable((*inhigh*) EN_cosq_val_in_dqPE5) ;
    method cosq_val_in_dqPE6(cosq_val_in_dqPE6) enable((*inhigh*) EN_cosq_val_in_dqPE6) ;
    method cosq_val_in_dqPE7(cosq_val_in_dqPE7) enable((*inhigh*) EN_cosq_val_in_dqPE7) ;
    method cosq_val_in_dqdPE1(cosq_val_in_dqdPE1) enable((*inhigh*) EN_cosq_val_in_dqdPE1) ;
    method cosq_val_in_dqdPE2(cosq_val_in_dqdPE2) enable((*inhigh*) EN_cosq_val_in_dqdPE2) ;
    method cosq_val_in_dqdPE3(cosq_val_in_dqdPE3) enable((*inhigh*) EN_cosq_val_in_dqdPE3) ;
    method cosq_val_in_dqdPE4(cosq_val_in_dqdPE4) enable((*inhigh*) EN_cosq_val_in_dqdPE4) ;
    method cosq_val_in_dqdPE5(cosq_val_in_dqdPE5) enable((*inhigh*) EN_cosq_val_in_dqdPE5) ;
    method cosq_val_in_dqdPE6(cosq_val_in_dqdPE6) enable((*inhigh*) EN_cosq_val_in_dqdPE6) ;
    method cosq_val_in_dqdPE7(cosq_val_in_dqdPE7) enable((*inhigh*) EN_cosq_val_in_dqdPE7) ;
    method qd_val_in_dqPE1(qd_val_in_dqPE1) enable((*inhigh*) EN_qd_val_in_dqPE1) ;
    method qd_val_in_dqPE2(qd_val_in_dqPE2) enable((*inhigh*) EN_qd_val_in_dqPE2) ;
    method qd_val_in_dqPE3(qd_val_in_dqPE3) enable((*inhigh*) EN_qd_val_in_dqPE3) ;
    method qd_val_in_dqPE4(qd_val_in_dqPE4) enable((*inhigh*) EN_qd_val_in_dqPE4) ;
    method qd_val_in_dqPE5(qd_val_in_dqPE5) enable((*inhigh*) EN_qd_val_in_dqPE5) ;
    method qd_val_in_dqPE6(qd_val_in_dqPE6) enable((*inhigh*) EN_qd_val_in_dqPE6) ;
    method qd_val_in_dqPE7(qd_val_in_dqPE7) enable((*inhigh*) EN_qd_val_in_dqPE7) ;
    method qd_val_in_dqdPE1(qd_val_in_dqdPE1) enable((*inhigh*) EN_qd_val_in_dqdPE1) ;
    method qd_val_in_dqdPE2(qd_val_in_dqdPE2) enable((*inhigh*) EN_qd_val_in_dqdPE2) ;
    method qd_val_in_dqdPE3(qd_val_in_dqdPE3) enable((*inhigh*) EN_qd_val_in_dqdPE3) ;
    method qd_val_in_dqdPE4(qd_val_in_dqdPE4) enable((*inhigh*) EN_qd_val_in_dqdPE4) ;
    method qd_val_in_dqdPE5(qd_val_in_dqdPE5) enable((*inhigh*) EN_qd_val_in_dqdPE5) ;
    method qd_val_in_dqdPE6(qd_val_in_dqdPE6) enable((*inhigh*) EN_qd_val_in_dqdPE6) ;
    method qd_val_in_dqdPE7(qd_val_in_dqdPE7) enable((*inhigh*) EN_qd_val_in_dqdPE7) ;

    method v_curr_vec_in_AX_dqPE1(v_curr_vec_in_AX_dqPE1) enable((*inhigh*) EN_v_curr_vec_in_AX_dqPE1) ;
    method v_curr_vec_in_AY_dqPE1(v_curr_vec_in_AY_dqPE1) enable((*inhigh*) EN_v_curr_vec_in_AY_dqPE1) ;
    method v_curr_vec_in_AZ_dqPE1(v_curr_vec_in_AZ_dqPE1) enable((*inhigh*) EN_v_curr_vec_in_AZ_dqPE1) ;
    method v_curr_vec_in_LX_dqPE1(v_curr_vec_in_LX_dqPE1) enable((*inhigh*) EN_v_curr_vec_in_LX_dqPE1) ;
    method v_curr_vec_in_LY_dqPE1(v_curr_vec_in_LY_dqPE1) enable((*inhigh*) EN_v_curr_vec_in_LY_dqPE1) ;
    method v_curr_vec_in_LZ_dqPE1(v_curr_vec_in_LZ_dqPE1) enable((*inhigh*) EN_v_curr_vec_in_LZ_dqPE1) ;
    method v_curr_vec_in_AX_dqPE2(v_curr_vec_in_AX_dqPE2) enable((*inhigh*) EN_v_curr_vec_in_AX_dqPE2) ;
    method v_curr_vec_in_AY_dqPE2(v_curr_vec_in_AY_dqPE2) enable((*inhigh*) EN_v_curr_vec_in_AY_dqPE2) ;
    method v_curr_vec_in_AZ_dqPE2(v_curr_vec_in_AZ_dqPE2) enable((*inhigh*) EN_v_curr_vec_in_AZ_dqPE2) ;
    method v_curr_vec_in_LX_dqPE2(v_curr_vec_in_LX_dqPE2) enable((*inhigh*) EN_v_curr_vec_in_LX_dqPE2) ;
    method v_curr_vec_in_LY_dqPE2(v_curr_vec_in_LY_dqPE2) enable((*inhigh*) EN_v_curr_vec_in_LY_dqPE2) ;
    method v_curr_vec_in_LZ_dqPE2(v_curr_vec_in_LZ_dqPE2) enable((*inhigh*) EN_v_curr_vec_in_LZ_dqPE2) ;
    method v_curr_vec_in_AX_dqPE3(v_curr_vec_in_AX_dqPE3) enable((*inhigh*) EN_v_curr_vec_in_AX_dqPE3) ;
    method v_curr_vec_in_AY_dqPE3(v_curr_vec_in_AY_dqPE3) enable((*inhigh*) EN_v_curr_vec_in_AY_dqPE3) ;
    method v_curr_vec_in_AZ_dqPE3(v_curr_vec_in_AZ_dqPE3) enable((*inhigh*) EN_v_curr_vec_in_AZ_dqPE3) ;
    method v_curr_vec_in_LX_dqPE3(v_curr_vec_in_LX_dqPE3) enable((*inhigh*) EN_v_curr_vec_in_LX_dqPE3) ;
    method v_curr_vec_in_LY_dqPE3(v_curr_vec_in_LY_dqPE3) enable((*inhigh*) EN_v_curr_vec_in_LY_dqPE3) ;
    method v_curr_vec_in_LZ_dqPE3(v_curr_vec_in_LZ_dqPE3) enable((*inhigh*) EN_v_curr_vec_in_LZ_dqPE3) ;
    method v_curr_vec_in_AX_dqPE4(v_curr_vec_in_AX_dqPE4) enable((*inhigh*) EN_v_curr_vec_in_AX_dqPE4) ;
    method v_curr_vec_in_AY_dqPE4(v_curr_vec_in_AY_dqPE4) enable((*inhigh*) EN_v_curr_vec_in_AY_dqPE4) ;
    method v_curr_vec_in_AZ_dqPE4(v_curr_vec_in_AZ_dqPE4) enable((*inhigh*) EN_v_curr_vec_in_AZ_dqPE4) ;
    method v_curr_vec_in_LX_dqPE4(v_curr_vec_in_LX_dqPE4) enable((*inhigh*) EN_v_curr_vec_in_LX_dqPE4) ;
    method v_curr_vec_in_LY_dqPE4(v_curr_vec_in_LY_dqPE4) enable((*inhigh*) EN_v_curr_vec_in_LY_dqPE4) ;
    method v_curr_vec_in_LZ_dqPE4(v_curr_vec_in_LZ_dqPE4) enable((*inhigh*) EN_v_curr_vec_in_LZ_dqPE4) ;
    method v_curr_vec_in_AX_dqPE5(v_curr_vec_in_AX_dqPE5) enable((*inhigh*) EN_v_curr_vec_in_AX_dqPE5) ;
    method v_curr_vec_in_AY_dqPE5(v_curr_vec_in_AY_dqPE5) enable((*inhigh*) EN_v_curr_vec_in_AY_dqPE5) ;
    method v_curr_vec_in_AZ_dqPE5(v_curr_vec_in_AZ_dqPE5) enable((*inhigh*) EN_v_curr_vec_in_AZ_dqPE5) ;
    method v_curr_vec_in_LX_dqPE5(v_curr_vec_in_LX_dqPE5) enable((*inhigh*) EN_v_curr_vec_in_LX_dqPE5) ;
    method v_curr_vec_in_LY_dqPE5(v_curr_vec_in_LY_dqPE5) enable((*inhigh*) EN_v_curr_vec_in_LY_dqPE5) ;
    method v_curr_vec_in_LZ_dqPE5(v_curr_vec_in_LZ_dqPE5) enable((*inhigh*) EN_v_curr_vec_in_LZ_dqPE5) ;
    method v_curr_vec_in_AX_dqPE6(v_curr_vec_in_AX_dqPE6) enable((*inhigh*) EN_v_curr_vec_in_AX_dqPE6) ;
    method v_curr_vec_in_AY_dqPE6(v_curr_vec_in_AY_dqPE6) enable((*inhigh*) EN_v_curr_vec_in_AY_dqPE6) ;
    method v_curr_vec_in_AZ_dqPE6(v_curr_vec_in_AZ_dqPE6) enable((*inhigh*) EN_v_curr_vec_in_AZ_dqPE6) ;
    method v_curr_vec_in_LX_dqPE6(v_curr_vec_in_LX_dqPE6) enable((*inhigh*) EN_v_curr_vec_in_LX_dqPE6) ;
    method v_curr_vec_in_LY_dqPE6(v_curr_vec_in_LY_dqPE6) enable((*inhigh*) EN_v_curr_vec_in_LY_dqPE6) ;
    method v_curr_vec_in_LZ_dqPE6(v_curr_vec_in_LZ_dqPE6) enable((*inhigh*) EN_v_curr_vec_in_LZ_dqPE6) ;
    method v_curr_vec_in_AX_dqPE7(v_curr_vec_in_AX_dqPE7) enable((*inhigh*) EN_v_curr_vec_in_AX_dqPE7) ;
    method v_curr_vec_in_AY_dqPE7(v_curr_vec_in_AY_dqPE7) enable((*inhigh*) EN_v_curr_vec_in_AY_dqPE7) ;
    method v_curr_vec_in_AZ_dqPE7(v_curr_vec_in_AZ_dqPE7) enable((*inhigh*) EN_v_curr_vec_in_AZ_dqPE7) ;
    method v_curr_vec_in_LX_dqPE7(v_curr_vec_in_LX_dqPE7) enable((*inhigh*) EN_v_curr_vec_in_LX_dqPE7) ;
    method v_curr_vec_in_LY_dqPE7(v_curr_vec_in_LY_dqPE7) enable((*inhigh*) EN_v_curr_vec_in_LY_dqPE7) ;
    method v_curr_vec_in_LZ_dqPE7(v_curr_vec_in_LZ_dqPE7) enable((*inhigh*) EN_v_curr_vec_in_LZ_dqPE7) ;
    method v_curr_vec_in_AX_dqdPE1(v_curr_vec_in_AX_dqdPE1) enable((*inhigh*) EN_v_curr_vec_in_AX_dqdPE1) ;
    method v_curr_vec_in_AY_dqdPE1(v_curr_vec_in_AY_dqdPE1) enable((*inhigh*) EN_v_curr_vec_in_AY_dqdPE1) ;
    method v_curr_vec_in_AZ_dqdPE1(v_curr_vec_in_AZ_dqdPE1) enable((*inhigh*) EN_v_curr_vec_in_AZ_dqdPE1) ;
    method v_curr_vec_in_LX_dqdPE1(v_curr_vec_in_LX_dqdPE1) enable((*inhigh*) EN_v_curr_vec_in_LX_dqdPE1) ;
    method v_curr_vec_in_LY_dqdPE1(v_curr_vec_in_LY_dqdPE1) enable((*inhigh*) EN_v_curr_vec_in_LY_dqdPE1) ;
    method v_curr_vec_in_LZ_dqdPE1(v_curr_vec_in_LZ_dqdPE1) enable((*inhigh*) EN_v_curr_vec_in_LZ_dqdPE1) ;
    method v_curr_vec_in_AX_dqdPE2(v_curr_vec_in_AX_dqdPE2) enable((*inhigh*) EN_v_curr_vec_in_AX_dqdPE2) ;
    method v_curr_vec_in_AY_dqdPE2(v_curr_vec_in_AY_dqdPE2) enable((*inhigh*) EN_v_curr_vec_in_AY_dqdPE2) ;
    method v_curr_vec_in_AZ_dqdPE2(v_curr_vec_in_AZ_dqdPE2) enable((*inhigh*) EN_v_curr_vec_in_AZ_dqdPE2) ;
    method v_curr_vec_in_LX_dqdPE2(v_curr_vec_in_LX_dqdPE2) enable((*inhigh*) EN_v_curr_vec_in_LX_dqdPE2) ;
    method v_curr_vec_in_LY_dqdPE2(v_curr_vec_in_LY_dqdPE2) enable((*inhigh*) EN_v_curr_vec_in_LY_dqdPE2) ;
    method v_curr_vec_in_LZ_dqdPE2(v_curr_vec_in_LZ_dqdPE2) enable((*inhigh*) EN_v_curr_vec_in_LZ_dqdPE2) ;
    method v_curr_vec_in_AX_dqdPE3(v_curr_vec_in_AX_dqdPE3) enable((*inhigh*) EN_v_curr_vec_in_AX_dqdPE3) ;
    method v_curr_vec_in_AY_dqdPE3(v_curr_vec_in_AY_dqdPE3) enable((*inhigh*) EN_v_curr_vec_in_AY_dqdPE3) ;
    method v_curr_vec_in_AZ_dqdPE3(v_curr_vec_in_AZ_dqdPE3) enable((*inhigh*) EN_v_curr_vec_in_AZ_dqdPE3) ;
    method v_curr_vec_in_LX_dqdPE3(v_curr_vec_in_LX_dqdPE3) enable((*inhigh*) EN_v_curr_vec_in_LX_dqdPE3) ;
    method v_curr_vec_in_LY_dqdPE3(v_curr_vec_in_LY_dqdPE3) enable((*inhigh*) EN_v_curr_vec_in_LY_dqdPE3) ;
    method v_curr_vec_in_LZ_dqdPE3(v_curr_vec_in_LZ_dqdPE3) enable((*inhigh*) EN_v_curr_vec_in_LZ_dqdPE3) ;
    method v_curr_vec_in_AX_dqdPE4(v_curr_vec_in_AX_dqdPE4) enable((*inhigh*) EN_v_curr_vec_in_AX_dqdPE4) ;
    method v_curr_vec_in_AY_dqdPE4(v_curr_vec_in_AY_dqdPE4) enable((*inhigh*) EN_v_curr_vec_in_AY_dqdPE4) ;
    method v_curr_vec_in_AZ_dqdPE4(v_curr_vec_in_AZ_dqdPE4) enable((*inhigh*) EN_v_curr_vec_in_AZ_dqdPE4) ;
    method v_curr_vec_in_LX_dqdPE4(v_curr_vec_in_LX_dqdPE4) enable((*inhigh*) EN_v_curr_vec_in_LX_dqdPE4) ;
    method v_curr_vec_in_LY_dqdPE4(v_curr_vec_in_LY_dqdPE4) enable((*inhigh*) EN_v_curr_vec_in_LY_dqdPE4) ;
    method v_curr_vec_in_LZ_dqdPE4(v_curr_vec_in_LZ_dqdPE4) enable((*inhigh*) EN_v_curr_vec_in_LZ_dqdPE4) ;
    method v_curr_vec_in_AX_dqdPE5(v_curr_vec_in_AX_dqdPE5) enable((*inhigh*) EN_v_curr_vec_in_AX_dqdPE5) ;
    method v_curr_vec_in_AY_dqdPE5(v_curr_vec_in_AY_dqdPE5) enable((*inhigh*) EN_v_curr_vec_in_AY_dqdPE5) ;
    method v_curr_vec_in_AZ_dqdPE5(v_curr_vec_in_AZ_dqdPE5) enable((*inhigh*) EN_v_curr_vec_in_AZ_dqdPE5) ;
    method v_curr_vec_in_LX_dqdPE5(v_curr_vec_in_LX_dqdPE5) enable((*inhigh*) EN_v_curr_vec_in_LX_dqdPE5) ;
    method v_curr_vec_in_LY_dqdPE5(v_curr_vec_in_LY_dqdPE5) enable((*inhigh*) EN_v_curr_vec_in_LY_dqdPE5) ;
    method v_curr_vec_in_LZ_dqdPE5(v_curr_vec_in_LZ_dqdPE5) enable((*inhigh*) EN_v_curr_vec_in_LZ_dqdPE5) ;
    method v_curr_vec_in_AX_dqdPE6(v_curr_vec_in_AX_dqdPE6) enable((*inhigh*) EN_v_curr_vec_in_AX_dqdPE6) ;
    method v_curr_vec_in_AY_dqdPE6(v_curr_vec_in_AY_dqdPE6) enable((*inhigh*) EN_v_curr_vec_in_AY_dqdPE6) ;
    method v_curr_vec_in_AZ_dqdPE6(v_curr_vec_in_AZ_dqdPE6) enable((*inhigh*) EN_v_curr_vec_in_AZ_dqdPE6) ;
    method v_curr_vec_in_LX_dqdPE6(v_curr_vec_in_LX_dqdPE6) enable((*inhigh*) EN_v_curr_vec_in_LX_dqdPE6) ;
    method v_curr_vec_in_LY_dqdPE6(v_curr_vec_in_LY_dqdPE6) enable((*inhigh*) EN_v_curr_vec_in_LY_dqdPE6) ;
    method v_curr_vec_in_LZ_dqdPE6(v_curr_vec_in_LZ_dqdPE6) enable((*inhigh*) EN_v_curr_vec_in_LZ_dqdPE6) ;
    method v_curr_vec_in_AX_dqdPE7(v_curr_vec_in_AX_dqdPE7) enable((*inhigh*) EN_v_curr_vec_in_AX_dqdPE7) ;
    method v_curr_vec_in_AY_dqdPE7(v_curr_vec_in_AY_dqdPE7) enable((*inhigh*) EN_v_curr_vec_in_AY_dqdPE7) ;
    method v_curr_vec_in_AZ_dqdPE7(v_curr_vec_in_AZ_dqdPE7) enable((*inhigh*) EN_v_curr_vec_in_AZ_dqdPE7) ;
    method v_curr_vec_in_LX_dqdPE7(v_curr_vec_in_LX_dqdPE7) enable((*inhigh*) EN_v_curr_vec_in_LX_dqdPE7) ;
    method v_curr_vec_in_LY_dqdPE7(v_curr_vec_in_LY_dqdPE7) enable((*inhigh*) EN_v_curr_vec_in_LY_dqdPE7) ;
    method v_curr_vec_in_LZ_dqdPE7(v_curr_vec_in_LZ_dqdPE7) enable((*inhigh*) EN_v_curr_vec_in_LZ_dqdPE7) ;
    method a_curr_vec_in_AX_dqPE1(a_curr_vec_in_AX_dqPE1) enable((*inhigh*) EN_a_curr_vec_in_AX_dqPE1) ;
    method a_curr_vec_in_AY_dqPE1(a_curr_vec_in_AY_dqPE1) enable((*inhigh*) EN_a_curr_vec_in_AY_dqPE1) ;
    method a_curr_vec_in_AZ_dqPE1(a_curr_vec_in_AZ_dqPE1) enable((*inhigh*) EN_a_curr_vec_in_AZ_dqPE1) ;
    method a_curr_vec_in_LX_dqPE1(a_curr_vec_in_LX_dqPE1) enable((*inhigh*) EN_a_curr_vec_in_LX_dqPE1) ;
    method a_curr_vec_in_LY_dqPE1(a_curr_vec_in_LY_dqPE1) enable((*inhigh*) EN_a_curr_vec_in_LY_dqPE1) ;
    method a_curr_vec_in_LZ_dqPE1(a_curr_vec_in_LZ_dqPE1) enable((*inhigh*) EN_a_curr_vec_in_LZ_dqPE1) ;
    method a_curr_vec_in_AX_dqPE2(a_curr_vec_in_AX_dqPE2) enable((*inhigh*) EN_a_curr_vec_in_AX_dqPE2) ;
    method a_curr_vec_in_AY_dqPE2(a_curr_vec_in_AY_dqPE2) enable((*inhigh*) EN_a_curr_vec_in_AY_dqPE2) ;
    method a_curr_vec_in_AZ_dqPE2(a_curr_vec_in_AZ_dqPE2) enable((*inhigh*) EN_a_curr_vec_in_AZ_dqPE2) ;
    method a_curr_vec_in_LX_dqPE2(a_curr_vec_in_LX_dqPE2) enable((*inhigh*) EN_a_curr_vec_in_LX_dqPE2) ;
    method a_curr_vec_in_LY_dqPE2(a_curr_vec_in_LY_dqPE2) enable((*inhigh*) EN_a_curr_vec_in_LY_dqPE2) ;
    method a_curr_vec_in_LZ_dqPE2(a_curr_vec_in_LZ_dqPE2) enable((*inhigh*) EN_a_curr_vec_in_LZ_dqPE2) ;
    method a_curr_vec_in_AX_dqPE3(a_curr_vec_in_AX_dqPE3) enable((*inhigh*) EN_a_curr_vec_in_AX_dqPE3) ;
    method a_curr_vec_in_AY_dqPE3(a_curr_vec_in_AY_dqPE3) enable((*inhigh*) EN_a_curr_vec_in_AY_dqPE3) ;
    method a_curr_vec_in_AZ_dqPE3(a_curr_vec_in_AZ_dqPE3) enable((*inhigh*) EN_a_curr_vec_in_AZ_dqPE3) ;
    method a_curr_vec_in_LX_dqPE3(a_curr_vec_in_LX_dqPE3) enable((*inhigh*) EN_a_curr_vec_in_LX_dqPE3) ;
    method a_curr_vec_in_LY_dqPE3(a_curr_vec_in_LY_dqPE3) enable((*inhigh*) EN_a_curr_vec_in_LY_dqPE3) ;
    method a_curr_vec_in_LZ_dqPE3(a_curr_vec_in_LZ_dqPE3) enable((*inhigh*) EN_a_curr_vec_in_LZ_dqPE3) ;
    method a_curr_vec_in_AX_dqPE4(a_curr_vec_in_AX_dqPE4) enable((*inhigh*) EN_a_curr_vec_in_AX_dqPE4) ;
    method a_curr_vec_in_AY_dqPE4(a_curr_vec_in_AY_dqPE4) enable((*inhigh*) EN_a_curr_vec_in_AY_dqPE4) ;
    method a_curr_vec_in_AZ_dqPE4(a_curr_vec_in_AZ_dqPE4) enable((*inhigh*) EN_a_curr_vec_in_AZ_dqPE4) ;
    method a_curr_vec_in_LX_dqPE4(a_curr_vec_in_LX_dqPE4) enable((*inhigh*) EN_a_curr_vec_in_LX_dqPE4) ;
    method a_curr_vec_in_LY_dqPE4(a_curr_vec_in_LY_dqPE4) enable((*inhigh*) EN_a_curr_vec_in_LY_dqPE4) ;
    method a_curr_vec_in_LZ_dqPE4(a_curr_vec_in_LZ_dqPE4) enable((*inhigh*) EN_a_curr_vec_in_LZ_dqPE4) ;
    method a_curr_vec_in_AX_dqPE5(a_curr_vec_in_AX_dqPE5) enable((*inhigh*) EN_a_curr_vec_in_AX_dqPE5) ;
    method a_curr_vec_in_AY_dqPE5(a_curr_vec_in_AY_dqPE5) enable((*inhigh*) EN_a_curr_vec_in_AY_dqPE5) ;
    method a_curr_vec_in_AZ_dqPE5(a_curr_vec_in_AZ_dqPE5) enable((*inhigh*) EN_a_curr_vec_in_AZ_dqPE5) ;
    method a_curr_vec_in_LX_dqPE5(a_curr_vec_in_LX_dqPE5) enable((*inhigh*) EN_a_curr_vec_in_LX_dqPE5) ;
    method a_curr_vec_in_LY_dqPE5(a_curr_vec_in_LY_dqPE5) enable((*inhigh*) EN_a_curr_vec_in_LY_dqPE5) ;
    method a_curr_vec_in_LZ_dqPE5(a_curr_vec_in_LZ_dqPE5) enable((*inhigh*) EN_a_curr_vec_in_LZ_dqPE5) ;
    method a_curr_vec_in_AX_dqPE6(a_curr_vec_in_AX_dqPE6) enable((*inhigh*) EN_a_curr_vec_in_AX_dqPE6) ;
    method a_curr_vec_in_AY_dqPE6(a_curr_vec_in_AY_dqPE6) enable((*inhigh*) EN_a_curr_vec_in_AY_dqPE6) ;
    method a_curr_vec_in_AZ_dqPE6(a_curr_vec_in_AZ_dqPE6) enable((*inhigh*) EN_a_curr_vec_in_AZ_dqPE6) ;
    method a_curr_vec_in_LX_dqPE6(a_curr_vec_in_LX_dqPE6) enable((*inhigh*) EN_a_curr_vec_in_LX_dqPE6) ;
    method a_curr_vec_in_LY_dqPE6(a_curr_vec_in_LY_dqPE6) enable((*inhigh*) EN_a_curr_vec_in_LY_dqPE6) ;
    method a_curr_vec_in_LZ_dqPE6(a_curr_vec_in_LZ_dqPE6) enable((*inhigh*) EN_a_curr_vec_in_LZ_dqPE6) ;
    method a_curr_vec_in_AX_dqPE7(a_curr_vec_in_AX_dqPE7) enable((*inhigh*) EN_a_curr_vec_in_AX_dqPE7) ;
    method a_curr_vec_in_AY_dqPE7(a_curr_vec_in_AY_dqPE7) enable((*inhigh*) EN_a_curr_vec_in_AY_dqPE7) ;
    method a_curr_vec_in_AZ_dqPE7(a_curr_vec_in_AZ_dqPE7) enable((*inhigh*) EN_a_curr_vec_in_AZ_dqPE7) ;
    method a_curr_vec_in_LX_dqPE7(a_curr_vec_in_LX_dqPE7) enable((*inhigh*) EN_a_curr_vec_in_LX_dqPE7) ;
    method a_curr_vec_in_LY_dqPE7(a_curr_vec_in_LY_dqPE7) enable((*inhigh*) EN_a_curr_vec_in_LY_dqPE7) ;
    method a_curr_vec_in_LZ_dqPE7(a_curr_vec_in_LZ_dqPE7) enable((*inhigh*) EN_a_curr_vec_in_LZ_dqPE7) ;
    method a_curr_vec_in_AX_dqdPE1(a_curr_vec_in_AX_dqdPE1) enable((*inhigh*) EN_a_curr_vec_in_AX_dqdPE1) ;
    method a_curr_vec_in_AY_dqdPE1(a_curr_vec_in_AY_dqdPE1) enable((*inhigh*) EN_a_curr_vec_in_AY_dqdPE1) ;
    method a_curr_vec_in_AZ_dqdPE1(a_curr_vec_in_AZ_dqdPE1) enable((*inhigh*) EN_a_curr_vec_in_AZ_dqdPE1) ;
    method a_curr_vec_in_LX_dqdPE1(a_curr_vec_in_LX_dqdPE1) enable((*inhigh*) EN_a_curr_vec_in_LX_dqdPE1) ;
    method a_curr_vec_in_LY_dqdPE1(a_curr_vec_in_LY_dqdPE1) enable((*inhigh*) EN_a_curr_vec_in_LY_dqdPE1) ;
    method a_curr_vec_in_LZ_dqdPE1(a_curr_vec_in_LZ_dqdPE1) enable((*inhigh*) EN_a_curr_vec_in_LZ_dqdPE1) ;
    method a_curr_vec_in_AX_dqdPE2(a_curr_vec_in_AX_dqdPE2) enable((*inhigh*) EN_a_curr_vec_in_AX_dqdPE2) ;
    method a_curr_vec_in_AY_dqdPE2(a_curr_vec_in_AY_dqdPE2) enable((*inhigh*) EN_a_curr_vec_in_AY_dqdPE2) ;
    method a_curr_vec_in_AZ_dqdPE2(a_curr_vec_in_AZ_dqdPE2) enable((*inhigh*) EN_a_curr_vec_in_AZ_dqdPE2) ;
    method a_curr_vec_in_LX_dqdPE2(a_curr_vec_in_LX_dqdPE2) enable((*inhigh*) EN_a_curr_vec_in_LX_dqdPE2) ;
    method a_curr_vec_in_LY_dqdPE2(a_curr_vec_in_LY_dqdPE2) enable((*inhigh*) EN_a_curr_vec_in_LY_dqdPE2) ;
    method a_curr_vec_in_LZ_dqdPE2(a_curr_vec_in_LZ_dqdPE2) enable((*inhigh*) EN_a_curr_vec_in_LZ_dqdPE2) ;
    method a_curr_vec_in_AX_dqdPE3(a_curr_vec_in_AX_dqdPE3) enable((*inhigh*) EN_a_curr_vec_in_AX_dqdPE3) ;
    method a_curr_vec_in_AY_dqdPE3(a_curr_vec_in_AY_dqdPE3) enable((*inhigh*) EN_a_curr_vec_in_AY_dqdPE3) ;
    method a_curr_vec_in_AZ_dqdPE3(a_curr_vec_in_AZ_dqdPE3) enable((*inhigh*) EN_a_curr_vec_in_AZ_dqdPE3) ;
    method a_curr_vec_in_LX_dqdPE3(a_curr_vec_in_LX_dqdPE3) enable((*inhigh*) EN_a_curr_vec_in_LX_dqdPE3) ;
    method a_curr_vec_in_LY_dqdPE3(a_curr_vec_in_LY_dqdPE3) enable((*inhigh*) EN_a_curr_vec_in_LY_dqdPE3) ;
    method a_curr_vec_in_LZ_dqdPE3(a_curr_vec_in_LZ_dqdPE3) enable((*inhigh*) EN_a_curr_vec_in_LZ_dqdPE3) ;
    method a_curr_vec_in_AX_dqdPE4(a_curr_vec_in_AX_dqdPE4) enable((*inhigh*) EN_a_curr_vec_in_AX_dqdPE4) ;
    method a_curr_vec_in_AY_dqdPE4(a_curr_vec_in_AY_dqdPE4) enable((*inhigh*) EN_a_curr_vec_in_AY_dqdPE4) ;
    method a_curr_vec_in_AZ_dqdPE4(a_curr_vec_in_AZ_dqdPE4) enable((*inhigh*) EN_a_curr_vec_in_AZ_dqdPE4) ;
    method a_curr_vec_in_LX_dqdPE4(a_curr_vec_in_LX_dqdPE4) enable((*inhigh*) EN_a_curr_vec_in_LX_dqdPE4) ;
    method a_curr_vec_in_LY_dqdPE4(a_curr_vec_in_LY_dqdPE4) enable((*inhigh*) EN_a_curr_vec_in_LY_dqdPE4) ;
    method a_curr_vec_in_LZ_dqdPE4(a_curr_vec_in_LZ_dqdPE4) enable((*inhigh*) EN_a_curr_vec_in_LZ_dqdPE4) ;
    method a_curr_vec_in_AX_dqdPE5(a_curr_vec_in_AX_dqdPE5) enable((*inhigh*) EN_a_curr_vec_in_AX_dqdPE5) ;
    method a_curr_vec_in_AY_dqdPE5(a_curr_vec_in_AY_dqdPE5) enable((*inhigh*) EN_a_curr_vec_in_AY_dqdPE5) ;
    method a_curr_vec_in_AZ_dqdPE5(a_curr_vec_in_AZ_dqdPE5) enable((*inhigh*) EN_a_curr_vec_in_AZ_dqdPE5) ;
    method a_curr_vec_in_LX_dqdPE5(a_curr_vec_in_LX_dqdPE5) enable((*inhigh*) EN_a_curr_vec_in_LX_dqdPE5) ;
    method a_curr_vec_in_LY_dqdPE5(a_curr_vec_in_LY_dqdPE5) enable((*inhigh*) EN_a_curr_vec_in_LY_dqdPE5) ;
    method a_curr_vec_in_LZ_dqdPE5(a_curr_vec_in_LZ_dqdPE5) enable((*inhigh*) EN_a_curr_vec_in_LZ_dqdPE5) ;
    method a_curr_vec_in_AX_dqdPE6(a_curr_vec_in_AX_dqdPE6) enable((*inhigh*) EN_a_curr_vec_in_AX_dqdPE6) ;
    method a_curr_vec_in_AY_dqdPE6(a_curr_vec_in_AY_dqdPE6) enable((*inhigh*) EN_a_curr_vec_in_AY_dqdPE6) ;
    method a_curr_vec_in_AZ_dqdPE6(a_curr_vec_in_AZ_dqdPE6) enable((*inhigh*) EN_a_curr_vec_in_AZ_dqdPE6) ;
    method a_curr_vec_in_LX_dqdPE6(a_curr_vec_in_LX_dqdPE6) enable((*inhigh*) EN_a_curr_vec_in_LX_dqdPE6) ;
    method a_curr_vec_in_LY_dqdPE6(a_curr_vec_in_LY_dqdPE6) enable((*inhigh*) EN_a_curr_vec_in_LY_dqdPE6) ;
    method a_curr_vec_in_LZ_dqdPE6(a_curr_vec_in_LZ_dqdPE6) enable((*inhigh*) EN_a_curr_vec_in_LZ_dqdPE6) ;
    method a_curr_vec_in_AX_dqdPE7(a_curr_vec_in_AX_dqdPE7) enable((*inhigh*) EN_a_curr_vec_in_AX_dqdPE7) ;
    method a_curr_vec_in_AY_dqdPE7(a_curr_vec_in_AY_dqdPE7) enable((*inhigh*) EN_a_curr_vec_in_AY_dqdPE7) ;
    method a_curr_vec_in_AZ_dqdPE7(a_curr_vec_in_AZ_dqdPE7) enable((*inhigh*) EN_a_curr_vec_in_AZ_dqdPE7) ;
    method a_curr_vec_in_LX_dqdPE7(a_curr_vec_in_LX_dqdPE7) enable((*inhigh*) EN_a_curr_vec_in_LX_dqdPE7) ;
    method a_curr_vec_in_LY_dqdPE7(a_curr_vec_in_LY_dqdPE7) enable((*inhigh*) EN_a_curr_vec_in_LY_dqdPE7) ;
    method a_curr_vec_in_LZ_dqdPE7(a_curr_vec_in_LZ_dqdPE7) enable((*inhigh*) EN_a_curr_vec_in_LZ_dqdPE7) ;
    method v_prev_vec_in_AX_dqPE1(v_prev_vec_in_AX_dqPE1) enable((*inhigh*) EN_v_prev_vec_in_AX_dqPE1) ;
    method v_prev_vec_in_AY_dqPE1(v_prev_vec_in_AY_dqPE1) enable((*inhigh*) EN_v_prev_vec_in_AY_dqPE1) ;
    method v_prev_vec_in_AZ_dqPE1(v_prev_vec_in_AZ_dqPE1) enable((*inhigh*) EN_v_prev_vec_in_AZ_dqPE1) ;
    method v_prev_vec_in_LX_dqPE1(v_prev_vec_in_LX_dqPE1) enable((*inhigh*) EN_v_prev_vec_in_LX_dqPE1) ;
    method v_prev_vec_in_LY_dqPE1(v_prev_vec_in_LY_dqPE1) enable((*inhigh*) EN_v_prev_vec_in_LY_dqPE1) ;
    method v_prev_vec_in_LZ_dqPE1(v_prev_vec_in_LZ_dqPE1) enable((*inhigh*) EN_v_prev_vec_in_LZ_dqPE1) ;
    method v_prev_vec_in_AX_dqPE2(v_prev_vec_in_AX_dqPE2) enable((*inhigh*) EN_v_prev_vec_in_AX_dqPE2) ;
    method v_prev_vec_in_AY_dqPE2(v_prev_vec_in_AY_dqPE2) enable((*inhigh*) EN_v_prev_vec_in_AY_dqPE2) ;
    method v_prev_vec_in_AZ_dqPE2(v_prev_vec_in_AZ_dqPE2) enable((*inhigh*) EN_v_prev_vec_in_AZ_dqPE2) ;
    method v_prev_vec_in_LX_dqPE2(v_prev_vec_in_LX_dqPE2) enable((*inhigh*) EN_v_prev_vec_in_LX_dqPE2) ;
    method v_prev_vec_in_LY_dqPE2(v_prev_vec_in_LY_dqPE2) enable((*inhigh*) EN_v_prev_vec_in_LY_dqPE2) ;
    method v_prev_vec_in_LZ_dqPE2(v_prev_vec_in_LZ_dqPE2) enable((*inhigh*) EN_v_prev_vec_in_LZ_dqPE2) ;
    method v_prev_vec_in_AX_dqPE3(v_prev_vec_in_AX_dqPE3) enable((*inhigh*) EN_v_prev_vec_in_AX_dqPE3) ;
    method v_prev_vec_in_AY_dqPE3(v_prev_vec_in_AY_dqPE3) enable((*inhigh*) EN_v_prev_vec_in_AY_dqPE3) ;
    method v_prev_vec_in_AZ_dqPE3(v_prev_vec_in_AZ_dqPE3) enable((*inhigh*) EN_v_prev_vec_in_AZ_dqPE3) ;
    method v_prev_vec_in_LX_dqPE3(v_prev_vec_in_LX_dqPE3) enable((*inhigh*) EN_v_prev_vec_in_LX_dqPE3) ;
    method v_prev_vec_in_LY_dqPE3(v_prev_vec_in_LY_dqPE3) enable((*inhigh*) EN_v_prev_vec_in_LY_dqPE3) ;
    method v_prev_vec_in_LZ_dqPE3(v_prev_vec_in_LZ_dqPE3) enable((*inhigh*) EN_v_prev_vec_in_LZ_dqPE3) ;
    method v_prev_vec_in_AX_dqPE4(v_prev_vec_in_AX_dqPE4) enable((*inhigh*) EN_v_prev_vec_in_AX_dqPE4) ;
    method v_prev_vec_in_AY_dqPE4(v_prev_vec_in_AY_dqPE4) enable((*inhigh*) EN_v_prev_vec_in_AY_dqPE4) ;
    method v_prev_vec_in_AZ_dqPE4(v_prev_vec_in_AZ_dqPE4) enable((*inhigh*) EN_v_prev_vec_in_AZ_dqPE4) ;
    method v_prev_vec_in_LX_dqPE4(v_prev_vec_in_LX_dqPE4) enable((*inhigh*) EN_v_prev_vec_in_LX_dqPE4) ;
    method v_prev_vec_in_LY_dqPE4(v_prev_vec_in_LY_dqPE4) enable((*inhigh*) EN_v_prev_vec_in_LY_dqPE4) ;
    method v_prev_vec_in_LZ_dqPE4(v_prev_vec_in_LZ_dqPE4) enable((*inhigh*) EN_v_prev_vec_in_LZ_dqPE4) ;
    method v_prev_vec_in_AX_dqPE5(v_prev_vec_in_AX_dqPE5) enable((*inhigh*) EN_v_prev_vec_in_AX_dqPE5) ;
    method v_prev_vec_in_AY_dqPE5(v_prev_vec_in_AY_dqPE5) enable((*inhigh*) EN_v_prev_vec_in_AY_dqPE5) ;
    method v_prev_vec_in_AZ_dqPE5(v_prev_vec_in_AZ_dqPE5) enable((*inhigh*) EN_v_prev_vec_in_AZ_dqPE5) ;
    method v_prev_vec_in_LX_dqPE5(v_prev_vec_in_LX_dqPE5) enable((*inhigh*) EN_v_prev_vec_in_LX_dqPE5) ;
    method v_prev_vec_in_LY_dqPE5(v_prev_vec_in_LY_dqPE5) enable((*inhigh*) EN_v_prev_vec_in_LY_dqPE5) ;
    method v_prev_vec_in_LZ_dqPE5(v_prev_vec_in_LZ_dqPE5) enable((*inhigh*) EN_v_prev_vec_in_LZ_dqPE5) ;
    method v_prev_vec_in_AX_dqPE6(v_prev_vec_in_AX_dqPE6) enable((*inhigh*) EN_v_prev_vec_in_AX_dqPE6) ;
    method v_prev_vec_in_AY_dqPE6(v_prev_vec_in_AY_dqPE6) enable((*inhigh*) EN_v_prev_vec_in_AY_dqPE6) ;
    method v_prev_vec_in_AZ_dqPE6(v_prev_vec_in_AZ_dqPE6) enable((*inhigh*) EN_v_prev_vec_in_AZ_dqPE6) ;
    method v_prev_vec_in_LX_dqPE6(v_prev_vec_in_LX_dqPE6) enable((*inhigh*) EN_v_prev_vec_in_LX_dqPE6) ;
    method v_prev_vec_in_LY_dqPE6(v_prev_vec_in_LY_dqPE6) enable((*inhigh*) EN_v_prev_vec_in_LY_dqPE6) ;
    method v_prev_vec_in_LZ_dqPE6(v_prev_vec_in_LZ_dqPE6) enable((*inhigh*) EN_v_prev_vec_in_LZ_dqPE6) ;
    method v_prev_vec_in_AX_dqPE7(v_prev_vec_in_AX_dqPE7) enable((*inhigh*) EN_v_prev_vec_in_AX_dqPE7) ;
    method v_prev_vec_in_AY_dqPE7(v_prev_vec_in_AY_dqPE7) enable((*inhigh*) EN_v_prev_vec_in_AY_dqPE7) ;
    method v_prev_vec_in_AZ_dqPE7(v_prev_vec_in_AZ_dqPE7) enable((*inhigh*) EN_v_prev_vec_in_AZ_dqPE7) ;
    method v_prev_vec_in_LX_dqPE7(v_prev_vec_in_LX_dqPE7) enable((*inhigh*) EN_v_prev_vec_in_LX_dqPE7) ;
    method v_prev_vec_in_LY_dqPE7(v_prev_vec_in_LY_dqPE7) enable((*inhigh*) EN_v_prev_vec_in_LY_dqPE7) ;
    method v_prev_vec_in_LZ_dqPE7(v_prev_vec_in_LZ_dqPE7) enable((*inhigh*) EN_v_prev_vec_in_LZ_dqPE7) ;
    method a_prev_vec_in_AX_dqPE1(a_prev_vec_in_AX_dqPE1) enable((*inhigh*) EN_a_prev_vec_in_AX_dqPE1) ;
    method a_prev_vec_in_AY_dqPE1(a_prev_vec_in_AY_dqPE1) enable((*inhigh*) EN_a_prev_vec_in_AY_dqPE1) ;
    method a_prev_vec_in_AZ_dqPE1(a_prev_vec_in_AZ_dqPE1) enable((*inhigh*) EN_a_prev_vec_in_AZ_dqPE1) ;
    method a_prev_vec_in_LX_dqPE1(a_prev_vec_in_LX_dqPE1) enable((*inhigh*) EN_a_prev_vec_in_LX_dqPE1) ;
    method a_prev_vec_in_LY_dqPE1(a_prev_vec_in_LY_dqPE1) enable((*inhigh*) EN_a_prev_vec_in_LY_dqPE1) ;
    method a_prev_vec_in_LZ_dqPE1(a_prev_vec_in_LZ_dqPE1) enable((*inhigh*) EN_a_prev_vec_in_LZ_dqPE1) ;
    method a_prev_vec_in_AX_dqPE2(a_prev_vec_in_AX_dqPE2) enable((*inhigh*) EN_a_prev_vec_in_AX_dqPE2) ;
    method a_prev_vec_in_AY_dqPE2(a_prev_vec_in_AY_dqPE2) enable((*inhigh*) EN_a_prev_vec_in_AY_dqPE2) ;
    method a_prev_vec_in_AZ_dqPE2(a_prev_vec_in_AZ_dqPE2) enable((*inhigh*) EN_a_prev_vec_in_AZ_dqPE2) ;
    method a_prev_vec_in_LX_dqPE2(a_prev_vec_in_LX_dqPE2) enable((*inhigh*) EN_a_prev_vec_in_LX_dqPE2) ;
    method a_prev_vec_in_LY_dqPE2(a_prev_vec_in_LY_dqPE2) enable((*inhigh*) EN_a_prev_vec_in_LY_dqPE2) ;
    method a_prev_vec_in_LZ_dqPE2(a_prev_vec_in_LZ_dqPE2) enable((*inhigh*) EN_a_prev_vec_in_LZ_dqPE2) ;
    method a_prev_vec_in_AX_dqPE3(a_prev_vec_in_AX_dqPE3) enable((*inhigh*) EN_a_prev_vec_in_AX_dqPE3) ;
    method a_prev_vec_in_AY_dqPE3(a_prev_vec_in_AY_dqPE3) enable((*inhigh*) EN_a_prev_vec_in_AY_dqPE3) ;
    method a_prev_vec_in_AZ_dqPE3(a_prev_vec_in_AZ_dqPE3) enable((*inhigh*) EN_a_prev_vec_in_AZ_dqPE3) ;
    method a_prev_vec_in_LX_dqPE3(a_prev_vec_in_LX_dqPE3) enable((*inhigh*) EN_a_prev_vec_in_LX_dqPE3) ;
    method a_prev_vec_in_LY_dqPE3(a_prev_vec_in_LY_dqPE3) enable((*inhigh*) EN_a_prev_vec_in_LY_dqPE3) ;
    method a_prev_vec_in_LZ_dqPE3(a_prev_vec_in_LZ_dqPE3) enable((*inhigh*) EN_a_prev_vec_in_LZ_dqPE3) ;
    method a_prev_vec_in_AX_dqPE4(a_prev_vec_in_AX_dqPE4) enable((*inhigh*) EN_a_prev_vec_in_AX_dqPE4) ;
    method a_prev_vec_in_AY_dqPE4(a_prev_vec_in_AY_dqPE4) enable((*inhigh*) EN_a_prev_vec_in_AY_dqPE4) ;
    method a_prev_vec_in_AZ_dqPE4(a_prev_vec_in_AZ_dqPE4) enable((*inhigh*) EN_a_prev_vec_in_AZ_dqPE4) ;
    method a_prev_vec_in_LX_dqPE4(a_prev_vec_in_LX_dqPE4) enable((*inhigh*) EN_a_prev_vec_in_LX_dqPE4) ;
    method a_prev_vec_in_LY_dqPE4(a_prev_vec_in_LY_dqPE4) enable((*inhigh*) EN_a_prev_vec_in_LY_dqPE4) ;
    method a_prev_vec_in_LZ_dqPE4(a_prev_vec_in_LZ_dqPE4) enable((*inhigh*) EN_a_prev_vec_in_LZ_dqPE4) ;
    method a_prev_vec_in_AX_dqPE5(a_prev_vec_in_AX_dqPE5) enable((*inhigh*) EN_a_prev_vec_in_AX_dqPE5) ;
    method a_prev_vec_in_AY_dqPE5(a_prev_vec_in_AY_dqPE5) enable((*inhigh*) EN_a_prev_vec_in_AY_dqPE5) ;
    method a_prev_vec_in_AZ_dqPE5(a_prev_vec_in_AZ_dqPE5) enable((*inhigh*) EN_a_prev_vec_in_AZ_dqPE5) ;
    method a_prev_vec_in_LX_dqPE5(a_prev_vec_in_LX_dqPE5) enable((*inhigh*) EN_a_prev_vec_in_LX_dqPE5) ;
    method a_prev_vec_in_LY_dqPE5(a_prev_vec_in_LY_dqPE5) enable((*inhigh*) EN_a_prev_vec_in_LY_dqPE5) ;
    method a_prev_vec_in_LZ_dqPE5(a_prev_vec_in_LZ_dqPE5) enable((*inhigh*) EN_a_prev_vec_in_LZ_dqPE5) ;
    method a_prev_vec_in_AX_dqPE6(a_prev_vec_in_AX_dqPE6) enable((*inhigh*) EN_a_prev_vec_in_AX_dqPE6) ;
    method a_prev_vec_in_AY_dqPE6(a_prev_vec_in_AY_dqPE6) enable((*inhigh*) EN_a_prev_vec_in_AY_dqPE6) ;
    method a_prev_vec_in_AZ_dqPE6(a_prev_vec_in_AZ_dqPE6) enable((*inhigh*) EN_a_prev_vec_in_AZ_dqPE6) ;
    method a_prev_vec_in_LX_dqPE6(a_prev_vec_in_LX_dqPE6) enable((*inhigh*) EN_a_prev_vec_in_LX_dqPE6) ;
    method a_prev_vec_in_LY_dqPE6(a_prev_vec_in_LY_dqPE6) enable((*inhigh*) EN_a_prev_vec_in_LY_dqPE6) ;
    method a_prev_vec_in_LZ_dqPE6(a_prev_vec_in_LZ_dqPE6) enable((*inhigh*) EN_a_prev_vec_in_LZ_dqPE6) ;
    method a_prev_vec_in_AX_dqPE7(a_prev_vec_in_AX_dqPE7) enable((*inhigh*) EN_a_prev_vec_in_AX_dqPE7) ;
    method a_prev_vec_in_AY_dqPE7(a_prev_vec_in_AY_dqPE7) enable((*inhigh*) EN_a_prev_vec_in_AY_dqPE7) ;
    method a_prev_vec_in_AZ_dqPE7(a_prev_vec_in_AZ_dqPE7) enable((*inhigh*) EN_a_prev_vec_in_AZ_dqPE7) ;
    method a_prev_vec_in_LX_dqPE7(a_prev_vec_in_LX_dqPE7) enable((*inhigh*) EN_a_prev_vec_in_LX_dqPE7) ;
    method a_prev_vec_in_LY_dqPE7(a_prev_vec_in_LY_dqPE7) enable((*inhigh*) EN_a_prev_vec_in_LY_dqPE7) ;
    method a_prev_vec_in_LZ_dqPE7(a_prev_vec_in_LZ_dqPE7) enable((*inhigh*) EN_a_prev_vec_in_LZ_dqPE7) ;

    method dvdq_prev_vec_in_AX_dqPE1(dvdq_prev_vec_in_AX_dqPE1) enable((*inhigh*) EN_dvdq_prev_vec_in_AX_dqPE1) ;
    method dvdq_prev_vec_in_AY_dqPE1(dvdq_prev_vec_in_AY_dqPE1) enable((*inhigh*) EN_dvdq_prev_vec_in_AY_dqPE1) ;
    method dvdq_prev_vec_in_AZ_dqPE1(dvdq_prev_vec_in_AZ_dqPE1) enable((*inhigh*) EN_dvdq_prev_vec_in_AZ_dqPE1) ;
    method dvdq_prev_vec_in_LX_dqPE1(dvdq_prev_vec_in_LX_dqPE1) enable((*inhigh*) EN_dvdq_prev_vec_in_LX_dqPE1) ;
    method dvdq_prev_vec_in_LY_dqPE1(dvdq_prev_vec_in_LY_dqPE1) enable((*inhigh*) EN_dvdq_prev_vec_in_LY_dqPE1) ;
    method dvdq_prev_vec_in_LZ_dqPE1(dvdq_prev_vec_in_LZ_dqPE1) enable((*inhigh*) EN_dvdq_prev_vec_in_LZ_dqPE1) ;
    method dvdq_prev_vec_in_AX_dqPE2(dvdq_prev_vec_in_AX_dqPE2) enable((*inhigh*) EN_dvdq_prev_vec_in_AX_dqPE2) ;
    method dvdq_prev_vec_in_AY_dqPE2(dvdq_prev_vec_in_AY_dqPE2) enable((*inhigh*) EN_dvdq_prev_vec_in_AY_dqPE2) ;
    method dvdq_prev_vec_in_AZ_dqPE2(dvdq_prev_vec_in_AZ_dqPE2) enable((*inhigh*) EN_dvdq_prev_vec_in_AZ_dqPE2) ;
    method dvdq_prev_vec_in_LX_dqPE2(dvdq_prev_vec_in_LX_dqPE2) enable((*inhigh*) EN_dvdq_prev_vec_in_LX_dqPE2) ;
    method dvdq_prev_vec_in_LY_dqPE2(dvdq_prev_vec_in_LY_dqPE2) enable((*inhigh*) EN_dvdq_prev_vec_in_LY_dqPE2) ;
    method dvdq_prev_vec_in_LZ_dqPE2(dvdq_prev_vec_in_LZ_dqPE2) enable((*inhigh*) EN_dvdq_prev_vec_in_LZ_dqPE2) ;
    method dvdq_prev_vec_in_AX_dqPE3(dvdq_prev_vec_in_AX_dqPE3) enable((*inhigh*) EN_dvdq_prev_vec_in_AX_dqPE3) ;
    method dvdq_prev_vec_in_AY_dqPE3(dvdq_prev_vec_in_AY_dqPE3) enable((*inhigh*) EN_dvdq_prev_vec_in_AY_dqPE3) ;
    method dvdq_prev_vec_in_AZ_dqPE3(dvdq_prev_vec_in_AZ_dqPE3) enable((*inhigh*) EN_dvdq_prev_vec_in_AZ_dqPE3) ;
    method dvdq_prev_vec_in_LX_dqPE3(dvdq_prev_vec_in_LX_dqPE3) enable((*inhigh*) EN_dvdq_prev_vec_in_LX_dqPE3) ;
    method dvdq_prev_vec_in_LY_dqPE3(dvdq_prev_vec_in_LY_dqPE3) enable((*inhigh*) EN_dvdq_prev_vec_in_LY_dqPE3) ;
    method dvdq_prev_vec_in_LZ_dqPE3(dvdq_prev_vec_in_LZ_dqPE3) enable((*inhigh*) EN_dvdq_prev_vec_in_LZ_dqPE3) ;
    method dvdq_prev_vec_in_AX_dqPE4(dvdq_prev_vec_in_AX_dqPE4) enable((*inhigh*) EN_dvdq_prev_vec_in_AX_dqPE4) ;
    method dvdq_prev_vec_in_AY_dqPE4(dvdq_prev_vec_in_AY_dqPE4) enable((*inhigh*) EN_dvdq_prev_vec_in_AY_dqPE4) ;
    method dvdq_prev_vec_in_AZ_dqPE4(dvdq_prev_vec_in_AZ_dqPE4) enable((*inhigh*) EN_dvdq_prev_vec_in_AZ_dqPE4) ;
    method dvdq_prev_vec_in_LX_dqPE4(dvdq_prev_vec_in_LX_dqPE4) enable((*inhigh*) EN_dvdq_prev_vec_in_LX_dqPE4) ;
    method dvdq_prev_vec_in_LY_dqPE4(dvdq_prev_vec_in_LY_dqPE4) enable((*inhigh*) EN_dvdq_prev_vec_in_LY_dqPE4) ;
    method dvdq_prev_vec_in_LZ_dqPE4(dvdq_prev_vec_in_LZ_dqPE4) enable((*inhigh*) EN_dvdq_prev_vec_in_LZ_dqPE4) ;
    method dvdq_prev_vec_in_AX_dqPE5(dvdq_prev_vec_in_AX_dqPE5) enable((*inhigh*) EN_dvdq_prev_vec_in_AX_dqPE5) ;
    method dvdq_prev_vec_in_AY_dqPE5(dvdq_prev_vec_in_AY_dqPE5) enable((*inhigh*) EN_dvdq_prev_vec_in_AY_dqPE5) ;
    method dvdq_prev_vec_in_AZ_dqPE5(dvdq_prev_vec_in_AZ_dqPE5) enable((*inhigh*) EN_dvdq_prev_vec_in_AZ_dqPE5) ;
    method dvdq_prev_vec_in_LX_dqPE5(dvdq_prev_vec_in_LX_dqPE5) enable((*inhigh*) EN_dvdq_prev_vec_in_LX_dqPE5) ;
    method dvdq_prev_vec_in_LY_dqPE5(dvdq_prev_vec_in_LY_dqPE5) enable((*inhigh*) EN_dvdq_prev_vec_in_LY_dqPE5) ;
    method dvdq_prev_vec_in_LZ_dqPE5(dvdq_prev_vec_in_LZ_dqPE5) enable((*inhigh*) EN_dvdq_prev_vec_in_LZ_dqPE5) ;
    method dvdq_prev_vec_in_AX_dqPE6(dvdq_prev_vec_in_AX_dqPE6) enable((*inhigh*) EN_dvdq_prev_vec_in_AX_dqPE6) ;
    method dvdq_prev_vec_in_AY_dqPE6(dvdq_prev_vec_in_AY_dqPE6) enable((*inhigh*) EN_dvdq_prev_vec_in_AY_dqPE6) ;
    method dvdq_prev_vec_in_AZ_dqPE6(dvdq_prev_vec_in_AZ_dqPE6) enable((*inhigh*) EN_dvdq_prev_vec_in_AZ_dqPE6) ;
    method dvdq_prev_vec_in_LX_dqPE6(dvdq_prev_vec_in_LX_dqPE6) enable((*inhigh*) EN_dvdq_prev_vec_in_LX_dqPE6) ;
    method dvdq_prev_vec_in_LY_dqPE6(dvdq_prev_vec_in_LY_dqPE6) enable((*inhigh*) EN_dvdq_prev_vec_in_LY_dqPE6) ;
    method dvdq_prev_vec_in_LZ_dqPE6(dvdq_prev_vec_in_LZ_dqPE6) enable((*inhigh*) EN_dvdq_prev_vec_in_LZ_dqPE6) ;
    method dvdq_prev_vec_in_AX_dqPE7(dvdq_prev_vec_in_AX_dqPE7) enable((*inhigh*) EN_dvdq_prev_vec_in_AX_dqPE7) ;
    method dvdq_prev_vec_in_AY_dqPE7(dvdq_prev_vec_in_AY_dqPE7) enable((*inhigh*) EN_dvdq_prev_vec_in_AY_dqPE7) ;
    method dvdq_prev_vec_in_AZ_dqPE7(dvdq_prev_vec_in_AZ_dqPE7) enable((*inhigh*) EN_dvdq_prev_vec_in_AZ_dqPE7) ;
    method dvdq_prev_vec_in_LX_dqPE7(dvdq_prev_vec_in_LX_dqPE7) enable((*inhigh*) EN_dvdq_prev_vec_in_LX_dqPE7) ;
    method dvdq_prev_vec_in_LY_dqPE7(dvdq_prev_vec_in_LY_dqPE7) enable((*inhigh*) EN_dvdq_prev_vec_in_LY_dqPE7) ;
    method dvdq_prev_vec_in_LZ_dqPE7(dvdq_prev_vec_in_LZ_dqPE7) enable((*inhigh*) EN_dvdq_prev_vec_in_LZ_dqPE7) ;
    method dvdqd_prev_vec_in_AX_dqdPE1(dvdqd_prev_vec_in_AX_dqdPE1) enable((*inhigh*) EN_dvdqd_prev_vec_in_AX_dqdPE1) ;
    method dvdqd_prev_vec_in_AY_dqdPE1(dvdqd_prev_vec_in_AY_dqdPE1) enable((*inhigh*) EN_dvdqd_prev_vec_in_AY_dqdPE1) ;
    method dvdqd_prev_vec_in_AZ_dqdPE1(dvdqd_prev_vec_in_AZ_dqdPE1) enable((*inhigh*) EN_dvdqd_prev_vec_in_AZ_dqdPE1) ;
    method dvdqd_prev_vec_in_LX_dqdPE1(dvdqd_prev_vec_in_LX_dqdPE1) enable((*inhigh*) EN_dvdqd_prev_vec_in_LX_dqdPE1) ;
    method dvdqd_prev_vec_in_LY_dqdPE1(dvdqd_prev_vec_in_LY_dqdPE1) enable((*inhigh*) EN_dvdqd_prev_vec_in_LY_dqdPE1) ;
    method dvdqd_prev_vec_in_LZ_dqdPE1(dvdqd_prev_vec_in_LZ_dqdPE1) enable((*inhigh*) EN_dvdqd_prev_vec_in_LZ_dqdPE1) ;
    method dvdqd_prev_vec_in_AX_dqdPE2(dvdqd_prev_vec_in_AX_dqdPE2) enable((*inhigh*) EN_dvdqd_prev_vec_in_AX_dqdPE2) ;
    method dvdqd_prev_vec_in_AY_dqdPE2(dvdqd_prev_vec_in_AY_dqdPE2) enable((*inhigh*) EN_dvdqd_prev_vec_in_AY_dqdPE2) ;
    method dvdqd_prev_vec_in_AZ_dqdPE2(dvdqd_prev_vec_in_AZ_dqdPE2) enable((*inhigh*) EN_dvdqd_prev_vec_in_AZ_dqdPE2) ;
    method dvdqd_prev_vec_in_LX_dqdPE2(dvdqd_prev_vec_in_LX_dqdPE2) enable((*inhigh*) EN_dvdqd_prev_vec_in_LX_dqdPE2) ;
    method dvdqd_prev_vec_in_LY_dqdPE2(dvdqd_prev_vec_in_LY_dqdPE2) enable((*inhigh*) EN_dvdqd_prev_vec_in_LY_dqdPE2) ;
    method dvdqd_prev_vec_in_LZ_dqdPE2(dvdqd_prev_vec_in_LZ_dqdPE2) enable((*inhigh*) EN_dvdqd_prev_vec_in_LZ_dqdPE2) ;
    method dvdqd_prev_vec_in_AX_dqdPE3(dvdqd_prev_vec_in_AX_dqdPE3) enable((*inhigh*) EN_dvdqd_prev_vec_in_AX_dqdPE3) ;
    method dvdqd_prev_vec_in_AY_dqdPE3(dvdqd_prev_vec_in_AY_dqdPE3) enable((*inhigh*) EN_dvdqd_prev_vec_in_AY_dqdPE3) ;
    method dvdqd_prev_vec_in_AZ_dqdPE3(dvdqd_prev_vec_in_AZ_dqdPE3) enable((*inhigh*) EN_dvdqd_prev_vec_in_AZ_dqdPE3) ;
    method dvdqd_prev_vec_in_LX_dqdPE3(dvdqd_prev_vec_in_LX_dqdPE3) enable((*inhigh*) EN_dvdqd_prev_vec_in_LX_dqdPE3) ;
    method dvdqd_prev_vec_in_LY_dqdPE3(dvdqd_prev_vec_in_LY_dqdPE3) enable((*inhigh*) EN_dvdqd_prev_vec_in_LY_dqdPE3) ;
    method dvdqd_prev_vec_in_LZ_dqdPE3(dvdqd_prev_vec_in_LZ_dqdPE3) enable((*inhigh*) EN_dvdqd_prev_vec_in_LZ_dqdPE3) ;
    method dvdqd_prev_vec_in_AX_dqdPE4(dvdqd_prev_vec_in_AX_dqdPE4) enable((*inhigh*) EN_dvdqd_prev_vec_in_AX_dqdPE4) ;
    method dvdqd_prev_vec_in_AY_dqdPE4(dvdqd_prev_vec_in_AY_dqdPE4) enable((*inhigh*) EN_dvdqd_prev_vec_in_AY_dqdPE4) ;
    method dvdqd_prev_vec_in_AZ_dqdPE4(dvdqd_prev_vec_in_AZ_dqdPE4) enable((*inhigh*) EN_dvdqd_prev_vec_in_AZ_dqdPE4) ;
    method dvdqd_prev_vec_in_LX_dqdPE4(dvdqd_prev_vec_in_LX_dqdPE4) enable((*inhigh*) EN_dvdqd_prev_vec_in_LX_dqdPE4) ;
    method dvdqd_prev_vec_in_LY_dqdPE4(dvdqd_prev_vec_in_LY_dqdPE4) enable((*inhigh*) EN_dvdqd_prev_vec_in_LY_dqdPE4) ;
    method dvdqd_prev_vec_in_LZ_dqdPE4(dvdqd_prev_vec_in_LZ_dqdPE4) enable((*inhigh*) EN_dvdqd_prev_vec_in_LZ_dqdPE4) ;
    method dvdqd_prev_vec_in_AX_dqdPE5(dvdqd_prev_vec_in_AX_dqdPE5) enable((*inhigh*) EN_dvdqd_prev_vec_in_AX_dqdPE5) ;
    method dvdqd_prev_vec_in_AY_dqdPE5(dvdqd_prev_vec_in_AY_dqdPE5) enable((*inhigh*) EN_dvdqd_prev_vec_in_AY_dqdPE5) ;
    method dvdqd_prev_vec_in_AZ_dqdPE5(dvdqd_prev_vec_in_AZ_dqdPE5) enable((*inhigh*) EN_dvdqd_prev_vec_in_AZ_dqdPE5) ;
    method dvdqd_prev_vec_in_LX_dqdPE5(dvdqd_prev_vec_in_LX_dqdPE5) enable((*inhigh*) EN_dvdqd_prev_vec_in_LX_dqdPE5) ;
    method dvdqd_prev_vec_in_LY_dqdPE5(dvdqd_prev_vec_in_LY_dqdPE5) enable((*inhigh*) EN_dvdqd_prev_vec_in_LY_dqdPE5) ;
    method dvdqd_prev_vec_in_LZ_dqdPE5(dvdqd_prev_vec_in_LZ_dqdPE5) enable((*inhigh*) EN_dvdqd_prev_vec_in_LZ_dqdPE5) ;
    method dvdqd_prev_vec_in_AX_dqdPE6(dvdqd_prev_vec_in_AX_dqdPE6) enable((*inhigh*) EN_dvdqd_prev_vec_in_AX_dqdPE6) ;
    method dvdqd_prev_vec_in_AY_dqdPE6(dvdqd_prev_vec_in_AY_dqdPE6) enable((*inhigh*) EN_dvdqd_prev_vec_in_AY_dqdPE6) ;
    method dvdqd_prev_vec_in_AZ_dqdPE6(dvdqd_prev_vec_in_AZ_dqdPE6) enable((*inhigh*) EN_dvdqd_prev_vec_in_AZ_dqdPE6) ;
    method dvdqd_prev_vec_in_LX_dqdPE6(dvdqd_prev_vec_in_LX_dqdPE6) enable((*inhigh*) EN_dvdqd_prev_vec_in_LX_dqdPE6) ;
    method dvdqd_prev_vec_in_LY_dqdPE6(dvdqd_prev_vec_in_LY_dqdPE6) enable((*inhigh*) EN_dvdqd_prev_vec_in_LY_dqdPE6) ;
    method dvdqd_prev_vec_in_LZ_dqdPE6(dvdqd_prev_vec_in_LZ_dqdPE6) enable((*inhigh*) EN_dvdqd_prev_vec_in_LZ_dqdPE6) ;
    method dvdqd_prev_vec_in_AX_dqdPE7(dvdqd_prev_vec_in_AX_dqdPE7) enable((*inhigh*) EN_dvdqd_prev_vec_in_AX_dqdPE7) ;
    method dvdqd_prev_vec_in_AY_dqdPE7(dvdqd_prev_vec_in_AY_dqdPE7) enable((*inhigh*) EN_dvdqd_prev_vec_in_AY_dqdPE7) ;
    method dvdqd_prev_vec_in_AZ_dqdPE7(dvdqd_prev_vec_in_AZ_dqdPE7) enable((*inhigh*) EN_dvdqd_prev_vec_in_AZ_dqdPE7) ;
    method dvdqd_prev_vec_in_LX_dqdPE7(dvdqd_prev_vec_in_LX_dqdPE7) enable((*inhigh*) EN_dvdqd_prev_vec_in_LX_dqdPE7) ;
    method dvdqd_prev_vec_in_LY_dqdPE7(dvdqd_prev_vec_in_LY_dqdPE7) enable((*inhigh*) EN_dvdqd_prev_vec_in_LY_dqdPE7) ;
    method dvdqd_prev_vec_in_LZ_dqdPE7(dvdqd_prev_vec_in_LZ_dqdPE7) enable((*inhigh*) EN_dvdqd_prev_vec_in_LZ_dqdPE7) ;
    method dadq_prev_vec_in_AX_dqPE1(dadq_prev_vec_in_AX_dqPE1) enable((*inhigh*) EN_dadq_prev_vec_in_AX_dqPE1) ;
    method dadq_prev_vec_in_AY_dqPE1(dadq_prev_vec_in_AY_dqPE1) enable((*inhigh*) EN_dadq_prev_vec_in_AY_dqPE1) ;
    method dadq_prev_vec_in_AZ_dqPE1(dadq_prev_vec_in_AZ_dqPE1) enable((*inhigh*) EN_dadq_prev_vec_in_AZ_dqPE1) ;
    method dadq_prev_vec_in_LX_dqPE1(dadq_prev_vec_in_LX_dqPE1) enable((*inhigh*) EN_dadq_prev_vec_in_LX_dqPE1) ;
    method dadq_prev_vec_in_LY_dqPE1(dadq_prev_vec_in_LY_dqPE1) enable((*inhigh*) EN_dadq_prev_vec_in_LY_dqPE1) ;
    method dadq_prev_vec_in_LZ_dqPE1(dadq_prev_vec_in_LZ_dqPE1) enable((*inhigh*) EN_dadq_prev_vec_in_LZ_dqPE1) ;
    method dadq_prev_vec_in_AX_dqPE2(dadq_prev_vec_in_AX_dqPE2) enable((*inhigh*) EN_dadq_prev_vec_in_AX_dqPE2) ;
    method dadq_prev_vec_in_AY_dqPE2(dadq_prev_vec_in_AY_dqPE2) enable((*inhigh*) EN_dadq_prev_vec_in_AY_dqPE2) ;
    method dadq_prev_vec_in_AZ_dqPE2(dadq_prev_vec_in_AZ_dqPE2) enable((*inhigh*) EN_dadq_prev_vec_in_AZ_dqPE2) ;
    method dadq_prev_vec_in_LX_dqPE2(dadq_prev_vec_in_LX_dqPE2) enable((*inhigh*) EN_dadq_prev_vec_in_LX_dqPE2) ;
    method dadq_prev_vec_in_LY_dqPE2(dadq_prev_vec_in_LY_dqPE2) enable((*inhigh*) EN_dadq_prev_vec_in_LY_dqPE2) ;
    method dadq_prev_vec_in_LZ_dqPE2(dadq_prev_vec_in_LZ_dqPE2) enable((*inhigh*) EN_dadq_prev_vec_in_LZ_dqPE2) ;
    method dadq_prev_vec_in_AX_dqPE3(dadq_prev_vec_in_AX_dqPE3) enable((*inhigh*) EN_dadq_prev_vec_in_AX_dqPE3) ;
    method dadq_prev_vec_in_AY_dqPE3(dadq_prev_vec_in_AY_dqPE3) enable((*inhigh*) EN_dadq_prev_vec_in_AY_dqPE3) ;
    method dadq_prev_vec_in_AZ_dqPE3(dadq_prev_vec_in_AZ_dqPE3) enable((*inhigh*) EN_dadq_prev_vec_in_AZ_dqPE3) ;
    method dadq_prev_vec_in_LX_dqPE3(dadq_prev_vec_in_LX_dqPE3) enable((*inhigh*) EN_dadq_prev_vec_in_LX_dqPE3) ;
    method dadq_prev_vec_in_LY_dqPE3(dadq_prev_vec_in_LY_dqPE3) enable((*inhigh*) EN_dadq_prev_vec_in_LY_dqPE3) ;
    method dadq_prev_vec_in_LZ_dqPE3(dadq_prev_vec_in_LZ_dqPE3) enable((*inhigh*) EN_dadq_prev_vec_in_LZ_dqPE3) ;
    method dadq_prev_vec_in_AX_dqPE4(dadq_prev_vec_in_AX_dqPE4) enable((*inhigh*) EN_dadq_prev_vec_in_AX_dqPE4) ;
    method dadq_prev_vec_in_AY_dqPE4(dadq_prev_vec_in_AY_dqPE4) enable((*inhigh*) EN_dadq_prev_vec_in_AY_dqPE4) ;
    method dadq_prev_vec_in_AZ_dqPE4(dadq_prev_vec_in_AZ_dqPE4) enable((*inhigh*) EN_dadq_prev_vec_in_AZ_dqPE4) ;
    method dadq_prev_vec_in_LX_dqPE4(dadq_prev_vec_in_LX_dqPE4) enable((*inhigh*) EN_dadq_prev_vec_in_LX_dqPE4) ;
    method dadq_prev_vec_in_LY_dqPE4(dadq_prev_vec_in_LY_dqPE4) enable((*inhigh*) EN_dadq_prev_vec_in_LY_dqPE4) ;
    method dadq_prev_vec_in_LZ_dqPE4(dadq_prev_vec_in_LZ_dqPE4) enable((*inhigh*) EN_dadq_prev_vec_in_LZ_dqPE4) ;
    method dadq_prev_vec_in_AX_dqPE5(dadq_prev_vec_in_AX_dqPE5) enable((*inhigh*) EN_dadq_prev_vec_in_AX_dqPE5) ;
    method dadq_prev_vec_in_AY_dqPE5(dadq_prev_vec_in_AY_dqPE5) enable((*inhigh*) EN_dadq_prev_vec_in_AY_dqPE5) ;
    method dadq_prev_vec_in_AZ_dqPE5(dadq_prev_vec_in_AZ_dqPE5) enable((*inhigh*) EN_dadq_prev_vec_in_AZ_dqPE5) ;
    method dadq_prev_vec_in_LX_dqPE5(dadq_prev_vec_in_LX_dqPE5) enable((*inhigh*) EN_dadq_prev_vec_in_LX_dqPE5) ;
    method dadq_prev_vec_in_LY_dqPE5(dadq_prev_vec_in_LY_dqPE5) enable((*inhigh*) EN_dadq_prev_vec_in_LY_dqPE5) ;
    method dadq_prev_vec_in_LZ_dqPE5(dadq_prev_vec_in_LZ_dqPE5) enable((*inhigh*) EN_dadq_prev_vec_in_LZ_dqPE5) ;
    method dadq_prev_vec_in_AX_dqPE6(dadq_prev_vec_in_AX_dqPE6) enable((*inhigh*) EN_dadq_prev_vec_in_AX_dqPE6) ;
    method dadq_prev_vec_in_AY_dqPE6(dadq_prev_vec_in_AY_dqPE6) enable((*inhigh*) EN_dadq_prev_vec_in_AY_dqPE6) ;
    method dadq_prev_vec_in_AZ_dqPE6(dadq_prev_vec_in_AZ_dqPE6) enable((*inhigh*) EN_dadq_prev_vec_in_AZ_dqPE6) ;
    method dadq_prev_vec_in_LX_dqPE6(dadq_prev_vec_in_LX_dqPE6) enable((*inhigh*) EN_dadq_prev_vec_in_LX_dqPE6) ;
    method dadq_prev_vec_in_LY_dqPE6(dadq_prev_vec_in_LY_dqPE6) enable((*inhigh*) EN_dadq_prev_vec_in_LY_dqPE6) ;
    method dadq_prev_vec_in_LZ_dqPE6(dadq_prev_vec_in_LZ_dqPE6) enable((*inhigh*) EN_dadq_prev_vec_in_LZ_dqPE6) ;
    method dadq_prev_vec_in_AX_dqPE7(dadq_prev_vec_in_AX_dqPE7) enable((*inhigh*) EN_dadq_prev_vec_in_AX_dqPE7) ;
    method dadq_prev_vec_in_AY_dqPE7(dadq_prev_vec_in_AY_dqPE7) enable((*inhigh*) EN_dadq_prev_vec_in_AY_dqPE7) ;
    method dadq_prev_vec_in_AZ_dqPE7(dadq_prev_vec_in_AZ_dqPE7) enable((*inhigh*) EN_dadq_prev_vec_in_AZ_dqPE7) ;
    method dadq_prev_vec_in_LX_dqPE7(dadq_prev_vec_in_LX_dqPE7) enable((*inhigh*) EN_dadq_prev_vec_in_LX_dqPE7) ;
    method dadq_prev_vec_in_LY_dqPE7(dadq_prev_vec_in_LY_dqPE7) enable((*inhigh*) EN_dadq_prev_vec_in_LY_dqPE7) ;
    method dadq_prev_vec_in_LZ_dqPE7(dadq_prev_vec_in_LZ_dqPE7) enable((*inhigh*) EN_dadq_prev_vec_in_LZ_dqPE7) ;
    method dadqd_prev_vec_in_AX_dqdPE1(dadqd_prev_vec_in_AX_dqdPE1) enable((*inhigh*) EN_dadqd_prev_vec_in_AX_dqdPE1) ;
    method dadqd_prev_vec_in_AY_dqdPE1(dadqd_prev_vec_in_AY_dqdPE1) enable((*inhigh*) EN_dadqd_prev_vec_in_AY_dqdPE1) ;
    method dadqd_prev_vec_in_AZ_dqdPE1(dadqd_prev_vec_in_AZ_dqdPE1) enable((*inhigh*) EN_dadqd_prev_vec_in_AZ_dqdPE1) ;
    method dadqd_prev_vec_in_LX_dqdPE1(dadqd_prev_vec_in_LX_dqdPE1) enable((*inhigh*) EN_dadqd_prev_vec_in_LX_dqdPE1) ;
    method dadqd_prev_vec_in_LY_dqdPE1(dadqd_prev_vec_in_LY_dqdPE1) enable((*inhigh*) EN_dadqd_prev_vec_in_LY_dqdPE1) ;
    method dadqd_prev_vec_in_LZ_dqdPE1(dadqd_prev_vec_in_LZ_dqdPE1) enable((*inhigh*) EN_dadqd_prev_vec_in_LZ_dqdPE1) ;
    method dadqd_prev_vec_in_AX_dqdPE2(dadqd_prev_vec_in_AX_dqdPE2) enable((*inhigh*) EN_dadqd_prev_vec_in_AX_dqdPE2) ;
    method dadqd_prev_vec_in_AY_dqdPE2(dadqd_prev_vec_in_AY_dqdPE2) enable((*inhigh*) EN_dadqd_prev_vec_in_AY_dqdPE2) ;
    method dadqd_prev_vec_in_AZ_dqdPE2(dadqd_prev_vec_in_AZ_dqdPE2) enable((*inhigh*) EN_dadqd_prev_vec_in_AZ_dqdPE2) ;
    method dadqd_prev_vec_in_LX_dqdPE2(dadqd_prev_vec_in_LX_dqdPE2) enable((*inhigh*) EN_dadqd_prev_vec_in_LX_dqdPE2) ;
    method dadqd_prev_vec_in_LY_dqdPE2(dadqd_prev_vec_in_LY_dqdPE2) enable((*inhigh*) EN_dadqd_prev_vec_in_LY_dqdPE2) ;
    method dadqd_prev_vec_in_LZ_dqdPE2(dadqd_prev_vec_in_LZ_dqdPE2) enable((*inhigh*) EN_dadqd_prev_vec_in_LZ_dqdPE2) ;
    method dadqd_prev_vec_in_AX_dqdPE3(dadqd_prev_vec_in_AX_dqdPE3) enable((*inhigh*) EN_dadqd_prev_vec_in_AX_dqdPE3) ;
    method dadqd_prev_vec_in_AY_dqdPE3(dadqd_prev_vec_in_AY_dqdPE3) enable((*inhigh*) EN_dadqd_prev_vec_in_AY_dqdPE3) ;
    method dadqd_prev_vec_in_AZ_dqdPE3(dadqd_prev_vec_in_AZ_dqdPE3) enable((*inhigh*) EN_dadqd_prev_vec_in_AZ_dqdPE3) ;
    method dadqd_prev_vec_in_LX_dqdPE3(dadqd_prev_vec_in_LX_dqdPE3) enable((*inhigh*) EN_dadqd_prev_vec_in_LX_dqdPE3) ;
    method dadqd_prev_vec_in_LY_dqdPE3(dadqd_prev_vec_in_LY_dqdPE3) enable((*inhigh*) EN_dadqd_prev_vec_in_LY_dqdPE3) ;
    method dadqd_prev_vec_in_LZ_dqdPE3(dadqd_prev_vec_in_LZ_dqdPE3) enable((*inhigh*) EN_dadqd_prev_vec_in_LZ_dqdPE3) ;
    method dadqd_prev_vec_in_AX_dqdPE4(dadqd_prev_vec_in_AX_dqdPE4) enable((*inhigh*) EN_dadqd_prev_vec_in_AX_dqdPE4) ;
    method dadqd_prev_vec_in_AY_dqdPE4(dadqd_prev_vec_in_AY_dqdPE4) enable((*inhigh*) EN_dadqd_prev_vec_in_AY_dqdPE4) ;
    method dadqd_prev_vec_in_AZ_dqdPE4(dadqd_prev_vec_in_AZ_dqdPE4) enable((*inhigh*) EN_dadqd_prev_vec_in_AZ_dqdPE4) ;
    method dadqd_prev_vec_in_LX_dqdPE4(dadqd_prev_vec_in_LX_dqdPE4) enable((*inhigh*) EN_dadqd_prev_vec_in_LX_dqdPE4) ;
    method dadqd_prev_vec_in_LY_dqdPE4(dadqd_prev_vec_in_LY_dqdPE4) enable((*inhigh*) EN_dadqd_prev_vec_in_LY_dqdPE4) ;
    method dadqd_prev_vec_in_LZ_dqdPE4(dadqd_prev_vec_in_LZ_dqdPE4) enable((*inhigh*) EN_dadqd_prev_vec_in_LZ_dqdPE4) ;
    method dadqd_prev_vec_in_AX_dqdPE5(dadqd_prev_vec_in_AX_dqdPE5) enable((*inhigh*) EN_dadqd_prev_vec_in_AX_dqdPE5) ;
    method dadqd_prev_vec_in_AY_dqdPE5(dadqd_prev_vec_in_AY_dqdPE5) enable((*inhigh*) EN_dadqd_prev_vec_in_AY_dqdPE5) ;
    method dadqd_prev_vec_in_AZ_dqdPE5(dadqd_prev_vec_in_AZ_dqdPE5) enable((*inhigh*) EN_dadqd_prev_vec_in_AZ_dqdPE5) ;
    method dadqd_prev_vec_in_LX_dqdPE5(dadqd_prev_vec_in_LX_dqdPE5) enable((*inhigh*) EN_dadqd_prev_vec_in_LX_dqdPE5) ;
    method dadqd_prev_vec_in_LY_dqdPE5(dadqd_prev_vec_in_LY_dqdPE5) enable((*inhigh*) EN_dadqd_prev_vec_in_LY_dqdPE5) ;
    method dadqd_prev_vec_in_LZ_dqdPE5(dadqd_prev_vec_in_LZ_dqdPE5) enable((*inhigh*) EN_dadqd_prev_vec_in_LZ_dqdPE5) ;
    method dadqd_prev_vec_in_AX_dqdPE6(dadqd_prev_vec_in_AX_dqdPE6) enable((*inhigh*) EN_dadqd_prev_vec_in_AX_dqdPE6) ;
    method dadqd_prev_vec_in_AY_dqdPE6(dadqd_prev_vec_in_AY_dqdPE6) enable((*inhigh*) EN_dadqd_prev_vec_in_AY_dqdPE6) ;
    method dadqd_prev_vec_in_AZ_dqdPE6(dadqd_prev_vec_in_AZ_dqdPE6) enable((*inhigh*) EN_dadqd_prev_vec_in_AZ_dqdPE6) ;
    method dadqd_prev_vec_in_LX_dqdPE6(dadqd_prev_vec_in_LX_dqdPE6) enable((*inhigh*) EN_dadqd_prev_vec_in_LX_dqdPE6) ;
    method dadqd_prev_vec_in_LY_dqdPE6(dadqd_prev_vec_in_LY_dqdPE6) enable((*inhigh*) EN_dadqd_prev_vec_in_LY_dqdPE6) ;
    method dadqd_prev_vec_in_LZ_dqdPE6(dadqd_prev_vec_in_LZ_dqdPE6) enable((*inhigh*) EN_dadqd_prev_vec_in_LZ_dqdPE6) ;
    method dadqd_prev_vec_in_AX_dqdPE7(dadqd_prev_vec_in_AX_dqdPE7) enable((*inhigh*) EN_dadqd_prev_vec_in_AX_dqdPE7) ;
    method dadqd_prev_vec_in_AY_dqdPE7(dadqd_prev_vec_in_AY_dqdPE7) enable((*inhigh*) EN_dadqd_prev_vec_in_AY_dqdPE7) ;
    method dadqd_prev_vec_in_AZ_dqdPE7(dadqd_prev_vec_in_AZ_dqdPE7) enable((*inhigh*) EN_dadqd_prev_vec_in_AZ_dqdPE7) ;
    method dadqd_prev_vec_in_LX_dqdPE7(dadqd_prev_vec_in_LX_dqdPE7) enable((*inhigh*) EN_dadqd_prev_vec_in_LX_dqdPE7) ;
    method dadqd_prev_vec_in_LY_dqdPE7(dadqd_prev_vec_in_LY_dqdPE7) enable((*inhigh*) EN_dadqd_prev_vec_in_LY_dqdPE7) ;
    method dadqd_prev_vec_in_LZ_dqdPE7(dadqd_prev_vec_in_LZ_dqdPE7) enable((*inhigh*) EN_dadqd_prev_vec_in_LZ_dqdPE7) ;

    method output_ready output_ready();

    method v_curr_vec_out_AX_rnea v_curr_vec_out_AX_rnea();
    method v_curr_vec_out_AY_rnea v_curr_vec_out_AY_rnea();
    method v_curr_vec_out_AZ_rnea v_curr_vec_out_AZ_rnea();
    method v_curr_vec_out_LX_rnea v_curr_vec_out_LX_rnea();
    method v_curr_vec_out_LY_rnea v_curr_vec_out_LY_rnea();
    method v_curr_vec_out_LZ_rnea v_curr_vec_out_LZ_rnea();
    method a_curr_vec_out_AX_rnea a_curr_vec_out_AX_rnea();
    method a_curr_vec_out_AY_rnea a_curr_vec_out_AY_rnea();
    method a_curr_vec_out_AZ_rnea a_curr_vec_out_AZ_rnea();
    method a_curr_vec_out_LX_rnea a_curr_vec_out_LX_rnea();
    method a_curr_vec_out_LY_rnea a_curr_vec_out_LY_rnea();
    method a_curr_vec_out_LZ_rnea a_curr_vec_out_LZ_rnea();
    method f_curr_vec_out_AX_rnea f_curr_vec_out_AX_rnea();
    method f_curr_vec_out_AY_rnea f_curr_vec_out_AY_rnea();
    method f_curr_vec_out_AZ_rnea f_curr_vec_out_AZ_rnea();
    method f_curr_vec_out_LX_rnea f_curr_vec_out_LX_rnea();
    method f_curr_vec_out_LY_rnea f_curr_vec_out_LY_rnea();
    method f_curr_vec_out_LZ_rnea f_curr_vec_out_LZ_rnea();

    method dfdq_curr_vec_out_AX_dqPE1 dfdq_curr_vec_out_AX_dqPE1();
    method dfdq_curr_vec_out_AY_dqPE1 dfdq_curr_vec_out_AY_dqPE1();
    method dfdq_curr_vec_out_AZ_dqPE1 dfdq_curr_vec_out_AZ_dqPE1();
    method dfdq_curr_vec_out_LX_dqPE1 dfdq_curr_vec_out_LX_dqPE1();
    method dfdq_curr_vec_out_LY_dqPE1 dfdq_curr_vec_out_LY_dqPE1();
    method dfdq_curr_vec_out_LZ_dqPE1 dfdq_curr_vec_out_LZ_dqPE1();
    method dfdq_curr_vec_out_AX_dqPE2 dfdq_curr_vec_out_AX_dqPE2();
    method dfdq_curr_vec_out_AY_dqPE2 dfdq_curr_vec_out_AY_dqPE2();
    method dfdq_curr_vec_out_AZ_dqPE2 dfdq_curr_vec_out_AZ_dqPE2();
    method dfdq_curr_vec_out_LX_dqPE2 dfdq_curr_vec_out_LX_dqPE2();
    method dfdq_curr_vec_out_LY_dqPE2 dfdq_curr_vec_out_LY_dqPE2();
    method dfdq_curr_vec_out_LZ_dqPE2 dfdq_curr_vec_out_LZ_dqPE2();
    method dfdq_curr_vec_out_AX_dqPE3 dfdq_curr_vec_out_AX_dqPE3();
    method dfdq_curr_vec_out_AY_dqPE3 dfdq_curr_vec_out_AY_dqPE3();
    method dfdq_curr_vec_out_AZ_dqPE3 dfdq_curr_vec_out_AZ_dqPE3();
    method dfdq_curr_vec_out_LX_dqPE3 dfdq_curr_vec_out_LX_dqPE3();
    method dfdq_curr_vec_out_LY_dqPE3 dfdq_curr_vec_out_LY_dqPE3();
    method dfdq_curr_vec_out_LZ_dqPE3 dfdq_curr_vec_out_LZ_dqPE3();
    method dfdq_curr_vec_out_AX_dqPE4 dfdq_curr_vec_out_AX_dqPE4();
    method dfdq_curr_vec_out_AY_dqPE4 dfdq_curr_vec_out_AY_dqPE4();
    method dfdq_curr_vec_out_AZ_dqPE4 dfdq_curr_vec_out_AZ_dqPE4();
    method dfdq_curr_vec_out_LX_dqPE4 dfdq_curr_vec_out_LX_dqPE4();
    method dfdq_curr_vec_out_LY_dqPE4 dfdq_curr_vec_out_LY_dqPE4();
    method dfdq_curr_vec_out_LZ_dqPE4 dfdq_curr_vec_out_LZ_dqPE4();
    method dfdq_curr_vec_out_AX_dqPE5 dfdq_curr_vec_out_AX_dqPE5();
    method dfdq_curr_vec_out_AY_dqPE5 dfdq_curr_vec_out_AY_dqPE5();
    method dfdq_curr_vec_out_AZ_dqPE5 dfdq_curr_vec_out_AZ_dqPE5();
    method dfdq_curr_vec_out_LX_dqPE5 dfdq_curr_vec_out_LX_dqPE5();
    method dfdq_curr_vec_out_LY_dqPE5 dfdq_curr_vec_out_LY_dqPE5();
    method dfdq_curr_vec_out_LZ_dqPE5 dfdq_curr_vec_out_LZ_dqPE5();
    method dfdq_curr_vec_out_AX_dqPE6 dfdq_curr_vec_out_AX_dqPE6();
    method dfdq_curr_vec_out_AY_dqPE6 dfdq_curr_vec_out_AY_dqPE6();
    method dfdq_curr_vec_out_AZ_dqPE6 dfdq_curr_vec_out_AZ_dqPE6();
    method dfdq_curr_vec_out_LX_dqPE6 dfdq_curr_vec_out_LX_dqPE6();
    method dfdq_curr_vec_out_LY_dqPE6 dfdq_curr_vec_out_LY_dqPE6();
    method dfdq_curr_vec_out_LZ_dqPE6 dfdq_curr_vec_out_LZ_dqPE6();
    method dfdq_curr_vec_out_AX_dqPE7 dfdq_curr_vec_out_AX_dqPE7();
    method dfdq_curr_vec_out_AY_dqPE7 dfdq_curr_vec_out_AY_dqPE7();
    method dfdq_curr_vec_out_AZ_dqPE7 dfdq_curr_vec_out_AZ_dqPE7();
    method dfdq_curr_vec_out_LX_dqPE7 dfdq_curr_vec_out_LX_dqPE7();
    method dfdq_curr_vec_out_LY_dqPE7 dfdq_curr_vec_out_LY_dqPE7();
    method dfdq_curr_vec_out_LZ_dqPE7 dfdq_curr_vec_out_LZ_dqPE7();
    method dfdqd_curr_vec_out_AX_dqdPE1 dfdqd_curr_vec_out_AX_dqdPE1();
    method dfdqd_curr_vec_out_AY_dqdPE1 dfdqd_curr_vec_out_AY_dqdPE1();
    method dfdqd_curr_vec_out_AZ_dqdPE1 dfdqd_curr_vec_out_AZ_dqdPE1();
    method dfdqd_curr_vec_out_LX_dqdPE1 dfdqd_curr_vec_out_LX_dqdPE1();
    method dfdqd_curr_vec_out_LY_dqdPE1 dfdqd_curr_vec_out_LY_dqdPE1();
    method dfdqd_curr_vec_out_LZ_dqdPE1 dfdqd_curr_vec_out_LZ_dqdPE1();
    method dfdqd_curr_vec_out_AX_dqdPE2 dfdqd_curr_vec_out_AX_dqdPE2();
    method dfdqd_curr_vec_out_AY_dqdPE2 dfdqd_curr_vec_out_AY_dqdPE2();
    method dfdqd_curr_vec_out_AZ_dqdPE2 dfdqd_curr_vec_out_AZ_dqdPE2();
    method dfdqd_curr_vec_out_LX_dqdPE2 dfdqd_curr_vec_out_LX_dqdPE2();
    method dfdqd_curr_vec_out_LY_dqdPE2 dfdqd_curr_vec_out_LY_dqdPE2();
    method dfdqd_curr_vec_out_LZ_dqdPE2 dfdqd_curr_vec_out_LZ_dqdPE2();
    method dfdqd_curr_vec_out_AX_dqdPE3 dfdqd_curr_vec_out_AX_dqdPE3();
    method dfdqd_curr_vec_out_AY_dqdPE3 dfdqd_curr_vec_out_AY_dqdPE3();
    method dfdqd_curr_vec_out_AZ_dqdPE3 dfdqd_curr_vec_out_AZ_dqdPE3();
    method dfdqd_curr_vec_out_LX_dqdPE3 dfdqd_curr_vec_out_LX_dqdPE3();
    method dfdqd_curr_vec_out_LY_dqdPE3 dfdqd_curr_vec_out_LY_dqdPE3();
    method dfdqd_curr_vec_out_LZ_dqdPE3 dfdqd_curr_vec_out_LZ_dqdPE3();
    method dfdqd_curr_vec_out_AX_dqdPE4 dfdqd_curr_vec_out_AX_dqdPE4();
    method dfdqd_curr_vec_out_AY_dqdPE4 dfdqd_curr_vec_out_AY_dqdPE4();
    method dfdqd_curr_vec_out_AZ_dqdPE4 dfdqd_curr_vec_out_AZ_dqdPE4();
    method dfdqd_curr_vec_out_LX_dqdPE4 dfdqd_curr_vec_out_LX_dqdPE4();
    method dfdqd_curr_vec_out_LY_dqdPE4 dfdqd_curr_vec_out_LY_dqdPE4();
    method dfdqd_curr_vec_out_LZ_dqdPE4 dfdqd_curr_vec_out_LZ_dqdPE4();
    method dfdqd_curr_vec_out_AX_dqdPE5 dfdqd_curr_vec_out_AX_dqdPE5();
    method dfdqd_curr_vec_out_AY_dqdPE5 dfdqd_curr_vec_out_AY_dqdPE5();
    method dfdqd_curr_vec_out_AZ_dqdPE5 dfdqd_curr_vec_out_AZ_dqdPE5();
    method dfdqd_curr_vec_out_LX_dqdPE5 dfdqd_curr_vec_out_LX_dqdPE5();
    method dfdqd_curr_vec_out_LY_dqdPE5 dfdqd_curr_vec_out_LY_dqdPE5();
    method dfdqd_curr_vec_out_LZ_dqdPE5 dfdqd_curr_vec_out_LZ_dqdPE5();
    method dfdqd_curr_vec_out_AX_dqdPE6 dfdqd_curr_vec_out_AX_dqdPE6();
    method dfdqd_curr_vec_out_AY_dqdPE6 dfdqd_curr_vec_out_AY_dqdPE6();
    method dfdqd_curr_vec_out_AZ_dqdPE6 dfdqd_curr_vec_out_AZ_dqdPE6();
    method dfdqd_curr_vec_out_LX_dqdPE6 dfdqd_curr_vec_out_LX_dqdPE6();
    method dfdqd_curr_vec_out_LY_dqdPE6 dfdqd_curr_vec_out_LY_dqdPE6();
    method dfdqd_curr_vec_out_LZ_dqdPE6 dfdqd_curr_vec_out_LZ_dqdPE6();
    method dfdqd_curr_vec_out_AX_dqdPE7 dfdqd_curr_vec_out_AX_dqdPE7();
    method dfdqd_curr_vec_out_AY_dqdPE7 dfdqd_curr_vec_out_AY_dqdPE7();
    method dfdqd_curr_vec_out_AZ_dqdPE7 dfdqd_curr_vec_out_AZ_dqdPE7();
    method dfdqd_curr_vec_out_LX_dqdPE7 dfdqd_curr_vec_out_LX_dqdPE7();
    method dfdqd_curr_vec_out_LY_dqdPE7 dfdqd_curr_vec_out_LY_dqdPE7();
    method dfdqd_curr_vec_out_LZ_dqdPE7 dfdqd_curr_vec_out_LZ_dqdPE7();

    method dvdq_curr_vec_out_AX_dqPE1 dvdq_curr_vec_out_AX_dqPE1();
    method dvdq_curr_vec_out_AY_dqPE1 dvdq_curr_vec_out_AY_dqPE1();
    method dvdq_curr_vec_out_AZ_dqPE1 dvdq_curr_vec_out_AZ_dqPE1();
    method dvdq_curr_vec_out_LX_dqPE1 dvdq_curr_vec_out_LX_dqPE1();
    method dvdq_curr_vec_out_LY_dqPE1 dvdq_curr_vec_out_LY_dqPE1();
    method dvdq_curr_vec_out_LZ_dqPE1 dvdq_curr_vec_out_LZ_dqPE1();
    method dvdq_curr_vec_out_AX_dqPE2 dvdq_curr_vec_out_AX_dqPE2();
    method dvdq_curr_vec_out_AY_dqPE2 dvdq_curr_vec_out_AY_dqPE2();
    method dvdq_curr_vec_out_AZ_dqPE2 dvdq_curr_vec_out_AZ_dqPE2();
    method dvdq_curr_vec_out_LX_dqPE2 dvdq_curr_vec_out_LX_dqPE2();
    method dvdq_curr_vec_out_LY_dqPE2 dvdq_curr_vec_out_LY_dqPE2();
    method dvdq_curr_vec_out_LZ_dqPE2 dvdq_curr_vec_out_LZ_dqPE2();
    method dvdq_curr_vec_out_AX_dqPE3 dvdq_curr_vec_out_AX_dqPE3();
    method dvdq_curr_vec_out_AY_dqPE3 dvdq_curr_vec_out_AY_dqPE3();
    method dvdq_curr_vec_out_AZ_dqPE3 dvdq_curr_vec_out_AZ_dqPE3();
    method dvdq_curr_vec_out_LX_dqPE3 dvdq_curr_vec_out_LX_dqPE3();
    method dvdq_curr_vec_out_LY_dqPE3 dvdq_curr_vec_out_LY_dqPE3();
    method dvdq_curr_vec_out_LZ_dqPE3 dvdq_curr_vec_out_LZ_dqPE3();
    method dvdq_curr_vec_out_AX_dqPE4 dvdq_curr_vec_out_AX_dqPE4();
    method dvdq_curr_vec_out_AY_dqPE4 dvdq_curr_vec_out_AY_dqPE4();
    method dvdq_curr_vec_out_AZ_dqPE4 dvdq_curr_vec_out_AZ_dqPE4();
    method dvdq_curr_vec_out_LX_dqPE4 dvdq_curr_vec_out_LX_dqPE4();
    method dvdq_curr_vec_out_LY_dqPE4 dvdq_curr_vec_out_LY_dqPE4();
    method dvdq_curr_vec_out_LZ_dqPE4 dvdq_curr_vec_out_LZ_dqPE4();
    method dvdq_curr_vec_out_AX_dqPE5 dvdq_curr_vec_out_AX_dqPE5();
    method dvdq_curr_vec_out_AY_dqPE5 dvdq_curr_vec_out_AY_dqPE5();
    method dvdq_curr_vec_out_AZ_dqPE5 dvdq_curr_vec_out_AZ_dqPE5();
    method dvdq_curr_vec_out_LX_dqPE5 dvdq_curr_vec_out_LX_dqPE5();
    method dvdq_curr_vec_out_LY_dqPE5 dvdq_curr_vec_out_LY_dqPE5();
    method dvdq_curr_vec_out_LZ_dqPE5 dvdq_curr_vec_out_LZ_dqPE5();
    method dvdq_curr_vec_out_AX_dqPE6 dvdq_curr_vec_out_AX_dqPE6();
    method dvdq_curr_vec_out_AY_dqPE6 dvdq_curr_vec_out_AY_dqPE6();
    method dvdq_curr_vec_out_AZ_dqPE6 dvdq_curr_vec_out_AZ_dqPE6();
    method dvdq_curr_vec_out_LX_dqPE6 dvdq_curr_vec_out_LX_dqPE6();
    method dvdq_curr_vec_out_LY_dqPE6 dvdq_curr_vec_out_LY_dqPE6();
    method dvdq_curr_vec_out_LZ_dqPE6 dvdq_curr_vec_out_LZ_dqPE6();
    method dvdq_curr_vec_out_AX_dqPE7 dvdq_curr_vec_out_AX_dqPE7();
    method dvdq_curr_vec_out_AY_dqPE7 dvdq_curr_vec_out_AY_dqPE7();
    method dvdq_curr_vec_out_AZ_dqPE7 dvdq_curr_vec_out_AZ_dqPE7();
    method dvdq_curr_vec_out_LX_dqPE7 dvdq_curr_vec_out_LX_dqPE7();
    method dvdq_curr_vec_out_LY_dqPE7 dvdq_curr_vec_out_LY_dqPE7();
    method dvdq_curr_vec_out_LZ_dqPE7 dvdq_curr_vec_out_LZ_dqPE7();
    method dvdqd_curr_vec_out_AX_dqdPE1 dvdqd_curr_vec_out_AX_dqdPE1();
    method dvdqd_curr_vec_out_AY_dqdPE1 dvdqd_curr_vec_out_AY_dqdPE1();
    method dvdqd_curr_vec_out_AZ_dqdPE1 dvdqd_curr_vec_out_AZ_dqdPE1();
    method dvdqd_curr_vec_out_LX_dqdPE1 dvdqd_curr_vec_out_LX_dqdPE1();
    method dvdqd_curr_vec_out_LY_dqdPE1 dvdqd_curr_vec_out_LY_dqdPE1();
    method dvdqd_curr_vec_out_LZ_dqdPE1 dvdqd_curr_vec_out_LZ_dqdPE1();
    method dvdqd_curr_vec_out_AX_dqdPE2 dvdqd_curr_vec_out_AX_dqdPE2();
    method dvdqd_curr_vec_out_AY_dqdPE2 dvdqd_curr_vec_out_AY_dqdPE2();
    method dvdqd_curr_vec_out_AZ_dqdPE2 dvdqd_curr_vec_out_AZ_dqdPE2();
    method dvdqd_curr_vec_out_LX_dqdPE2 dvdqd_curr_vec_out_LX_dqdPE2();
    method dvdqd_curr_vec_out_LY_dqdPE2 dvdqd_curr_vec_out_LY_dqdPE2();
    method dvdqd_curr_vec_out_LZ_dqdPE2 dvdqd_curr_vec_out_LZ_dqdPE2();
    method dvdqd_curr_vec_out_AX_dqdPE3 dvdqd_curr_vec_out_AX_dqdPE3();
    method dvdqd_curr_vec_out_AY_dqdPE3 dvdqd_curr_vec_out_AY_dqdPE3();
    method dvdqd_curr_vec_out_AZ_dqdPE3 dvdqd_curr_vec_out_AZ_dqdPE3();
    method dvdqd_curr_vec_out_LX_dqdPE3 dvdqd_curr_vec_out_LX_dqdPE3();
    method dvdqd_curr_vec_out_LY_dqdPE3 dvdqd_curr_vec_out_LY_dqdPE3();
    method dvdqd_curr_vec_out_LZ_dqdPE3 dvdqd_curr_vec_out_LZ_dqdPE3();
    method dvdqd_curr_vec_out_AX_dqdPE4 dvdqd_curr_vec_out_AX_dqdPE4();
    method dvdqd_curr_vec_out_AY_dqdPE4 dvdqd_curr_vec_out_AY_dqdPE4();
    method dvdqd_curr_vec_out_AZ_dqdPE4 dvdqd_curr_vec_out_AZ_dqdPE4();
    method dvdqd_curr_vec_out_LX_dqdPE4 dvdqd_curr_vec_out_LX_dqdPE4();
    method dvdqd_curr_vec_out_LY_dqdPE4 dvdqd_curr_vec_out_LY_dqdPE4();
    method dvdqd_curr_vec_out_LZ_dqdPE4 dvdqd_curr_vec_out_LZ_dqdPE4();
    method dvdqd_curr_vec_out_AX_dqdPE5 dvdqd_curr_vec_out_AX_dqdPE5();
    method dvdqd_curr_vec_out_AY_dqdPE5 dvdqd_curr_vec_out_AY_dqdPE5();
    method dvdqd_curr_vec_out_AZ_dqdPE5 dvdqd_curr_vec_out_AZ_dqdPE5();
    method dvdqd_curr_vec_out_LX_dqdPE5 dvdqd_curr_vec_out_LX_dqdPE5();
    method dvdqd_curr_vec_out_LY_dqdPE5 dvdqd_curr_vec_out_LY_dqdPE5();
    method dvdqd_curr_vec_out_LZ_dqdPE5 dvdqd_curr_vec_out_LZ_dqdPE5();
    method dvdqd_curr_vec_out_AX_dqdPE6 dvdqd_curr_vec_out_AX_dqdPE6();
    method dvdqd_curr_vec_out_AY_dqdPE6 dvdqd_curr_vec_out_AY_dqdPE6();
    method dvdqd_curr_vec_out_AZ_dqdPE6 dvdqd_curr_vec_out_AZ_dqdPE6();
    method dvdqd_curr_vec_out_LX_dqdPE6 dvdqd_curr_vec_out_LX_dqdPE6();
    method dvdqd_curr_vec_out_LY_dqdPE6 dvdqd_curr_vec_out_LY_dqdPE6();
    method dvdqd_curr_vec_out_LZ_dqdPE6 dvdqd_curr_vec_out_LZ_dqdPE6();
    method dvdqd_curr_vec_out_AX_dqdPE7 dvdqd_curr_vec_out_AX_dqdPE7();
    method dvdqd_curr_vec_out_AY_dqdPE7 dvdqd_curr_vec_out_AY_dqdPE7();
    method dvdqd_curr_vec_out_AZ_dqdPE7 dvdqd_curr_vec_out_AZ_dqdPE7();
    method dvdqd_curr_vec_out_LX_dqdPE7 dvdqd_curr_vec_out_LX_dqdPE7();
    method dvdqd_curr_vec_out_LY_dqdPE7 dvdqd_curr_vec_out_LY_dqdPE7();
    method dvdqd_curr_vec_out_LZ_dqdPE7 dvdqd_curr_vec_out_LZ_dqdPE7();
    method dadq_curr_vec_out_AX_dqPE1 dadq_curr_vec_out_AX_dqPE1();
    method dadq_curr_vec_out_AY_dqPE1 dadq_curr_vec_out_AY_dqPE1();
    method dadq_curr_vec_out_AZ_dqPE1 dadq_curr_vec_out_AZ_dqPE1();
    method dadq_curr_vec_out_LX_dqPE1 dadq_curr_vec_out_LX_dqPE1();
    method dadq_curr_vec_out_LY_dqPE1 dadq_curr_vec_out_LY_dqPE1();
    method dadq_curr_vec_out_LZ_dqPE1 dadq_curr_vec_out_LZ_dqPE1();
    method dadq_curr_vec_out_AX_dqPE2 dadq_curr_vec_out_AX_dqPE2();
    method dadq_curr_vec_out_AY_dqPE2 dadq_curr_vec_out_AY_dqPE2();
    method dadq_curr_vec_out_AZ_dqPE2 dadq_curr_vec_out_AZ_dqPE2();
    method dadq_curr_vec_out_LX_dqPE2 dadq_curr_vec_out_LX_dqPE2();
    method dadq_curr_vec_out_LY_dqPE2 dadq_curr_vec_out_LY_dqPE2();
    method dadq_curr_vec_out_LZ_dqPE2 dadq_curr_vec_out_LZ_dqPE2();
    method dadq_curr_vec_out_AX_dqPE3 dadq_curr_vec_out_AX_dqPE3();
    method dadq_curr_vec_out_AY_dqPE3 dadq_curr_vec_out_AY_dqPE3();
    method dadq_curr_vec_out_AZ_dqPE3 dadq_curr_vec_out_AZ_dqPE3();
    method dadq_curr_vec_out_LX_dqPE3 dadq_curr_vec_out_LX_dqPE3();
    method dadq_curr_vec_out_LY_dqPE3 dadq_curr_vec_out_LY_dqPE3();
    method dadq_curr_vec_out_LZ_dqPE3 dadq_curr_vec_out_LZ_dqPE3();
    method dadq_curr_vec_out_AX_dqPE4 dadq_curr_vec_out_AX_dqPE4();
    method dadq_curr_vec_out_AY_dqPE4 dadq_curr_vec_out_AY_dqPE4();
    method dadq_curr_vec_out_AZ_dqPE4 dadq_curr_vec_out_AZ_dqPE4();
    method dadq_curr_vec_out_LX_dqPE4 dadq_curr_vec_out_LX_dqPE4();
    method dadq_curr_vec_out_LY_dqPE4 dadq_curr_vec_out_LY_dqPE4();
    method dadq_curr_vec_out_LZ_dqPE4 dadq_curr_vec_out_LZ_dqPE4();
    method dadq_curr_vec_out_AX_dqPE5 dadq_curr_vec_out_AX_dqPE5();
    method dadq_curr_vec_out_AY_dqPE5 dadq_curr_vec_out_AY_dqPE5();
    method dadq_curr_vec_out_AZ_dqPE5 dadq_curr_vec_out_AZ_dqPE5();
    method dadq_curr_vec_out_LX_dqPE5 dadq_curr_vec_out_LX_dqPE5();
    method dadq_curr_vec_out_LY_dqPE5 dadq_curr_vec_out_LY_dqPE5();
    method dadq_curr_vec_out_LZ_dqPE5 dadq_curr_vec_out_LZ_dqPE5();
    method dadq_curr_vec_out_AX_dqPE6 dadq_curr_vec_out_AX_dqPE6();
    method dadq_curr_vec_out_AY_dqPE6 dadq_curr_vec_out_AY_dqPE6();
    method dadq_curr_vec_out_AZ_dqPE6 dadq_curr_vec_out_AZ_dqPE6();
    method dadq_curr_vec_out_LX_dqPE6 dadq_curr_vec_out_LX_dqPE6();
    method dadq_curr_vec_out_LY_dqPE6 dadq_curr_vec_out_LY_dqPE6();
    method dadq_curr_vec_out_LZ_dqPE6 dadq_curr_vec_out_LZ_dqPE6();
    method dadq_curr_vec_out_AX_dqPE7 dadq_curr_vec_out_AX_dqPE7();
    method dadq_curr_vec_out_AY_dqPE7 dadq_curr_vec_out_AY_dqPE7();
    method dadq_curr_vec_out_AZ_dqPE7 dadq_curr_vec_out_AZ_dqPE7();
    method dadq_curr_vec_out_LX_dqPE7 dadq_curr_vec_out_LX_dqPE7();
    method dadq_curr_vec_out_LY_dqPE7 dadq_curr_vec_out_LY_dqPE7();
    method dadq_curr_vec_out_LZ_dqPE7 dadq_curr_vec_out_LZ_dqPE7();
    method dadqd_curr_vec_out_AX_dqdPE1 dadqd_curr_vec_out_AX_dqdPE1();
    method dadqd_curr_vec_out_AY_dqdPE1 dadqd_curr_vec_out_AY_dqdPE1();
    method dadqd_curr_vec_out_AZ_dqdPE1 dadqd_curr_vec_out_AZ_dqdPE1();
    method dadqd_curr_vec_out_LX_dqdPE1 dadqd_curr_vec_out_LX_dqdPE1();
    method dadqd_curr_vec_out_LY_dqdPE1 dadqd_curr_vec_out_LY_dqdPE1();
    method dadqd_curr_vec_out_LZ_dqdPE1 dadqd_curr_vec_out_LZ_dqdPE1();
    method dadqd_curr_vec_out_AX_dqdPE2 dadqd_curr_vec_out_AX_dqdPE2();
    method dadqd_curr_vec_out_AY_dqdPE2 dadqd_curr_vec_out_AY_dqdPE2();
    method dadqd_curr_vec_out_AZ_dqdPE2 dadqd_curr_vec_out_AZ_dqdPE2();
    method dadqd_curr_vec_out_LX_dqdPE2 dadqd_curr_vec_out_LX_dqdPE2();
    method dadqd_curr_vec_out_LY_dqdPE2 dadqd_curr_vec_out_LY_dqdPE2();
    method dadqd_curr_vec_out_LZ_dqdPE2 dadqd_curr_vec_out_LZ_dqdPE2();
    method dadqd_curr_vec_out_AX_dqdPE3 dadqd_curr_vec_out_AX_dqdPE3();
    method dadqd_curr_vec_out_AY_dqdPE3 dadqd_curr_vec_out_AY_dqdPE3();
    method dadqd_curr_vec_out_AZ_dqdPE3 dadqd_curr_vec_out_AZ_dqdPE3();
    method dadqd_curr_vec_out_LX_dqdPE3 dadqd_curr_vec_out_LX_dqdPE3();
    method dadqd_curr_vec_out_LY_dqdPE3 dadqd_curr_vec_out_LY_dqdPE3();
    method dadqd_curr_vec_out_LZ_dqdPE3 dadqd_curr_vec_out_LZ_dqdPE3();
    method dadqd_curr_vec_out_AX_dqdPE4 dadqd_curr_vec_out_AX_dqdPE4();
    method dadqd_curr_vec_out_AY_dqdPE4 dadqd_curr_vec_out_AY_dqdPE4();
    method dadqd_curr_vec_out_AZ_dqdPE4 dadqd_curr_vec_out_AZ_dqdPE4();
    method dadqd_curr_vec_out_LX_dqdPE4 dadqd_curr_vec_out_LX_dqdPE4();
    method dadqd_curr_vec_out_LY_dqdPE4 dadqd_curr_vec_out_LY_dqdPE4();
    method dadqd_curr_vec_out_LZ_dqdPE4 dadqd_curr_vec_out_LZ_dqdPE4();
    method dadqd_curr_vec_out_AX_dqdPE5 dadqd_curr_vec_out_AX_dqdPE5();
    method dadqd_curr_vec_out_AY_dqdPE5 dadqd_curr_vec_out_AY_dqdPE5();
    method dadqd_curr_vec_out_AZ_dqdPE5 dadqd_curr_vec_out_AZ_dqdPE5();
    method dadqd_curr_vec_out_LX_dqdPE5 dadqd_curr_vec_out_LX_dqdPE5();
    method dadqd_curr_vec_out_LY_dqdPE5 dadqd_curr_vec_out_LY_dqdPE5();
    method dadqd_curr_vec_out_LZ_dqdPE5 dadqd_curr_vec_out_LZ_dqdPE5();
    method dadqd_curr_vec_out_AX_dqdPE6 dadqd_curr_vec_out_AX_dqdPE6();
    method dadqd_curr_vec_out_AY_dqdPE6 dadqd_curr_vec_out_AY_dqdPE6();
    method dadqd_curr_vec_out_AZ_dqdPE6 dadqd_curr_vec_out_AZ_dqdPE6();
    method dadqd_curr_vec_out_LX_dqdPE6 dadqd_curr_vec_out_LX_dqdPE6();
    method dadqd_curr_vec_out_LY_dqdPE6 dadqd_curr_vec_out_LY_dqdPE6();
    method dadqd_curr_vec_out_LZ_dqdPE6 dadqd_curr_vec_out_LZ_dqdPE6();
    method dadqd_curr_vec_out_AX_dqdPE7 dadqd_curr_vec_out_AX_dqdPE7();
    method dadqd_curr_vec_out_AY_dqdPE7 dadqd_curr_vec_out_AY_dqdPE7();
    method dadqd_curr_vec_out_AZ_dqdPE7 dadqd_curr_vec_out_AZ_dqdPE7();
    method dadqd_curr_vec_out_LX_dqdPE7 dadqd_curr_vec_out_LX_dqdPE7();
    method dadqd_curr_vec_out_LY_dqdPE7 dadqd_curr_vec_out_LY_dqdPE7();
    method dadqd_curr_vec_out_LZ_dqdPE7 dadqd_curr_vec_out_LZ_dqdPE7();

    schedule (
        get_data, link_in_rnea, sinq_val_in_rnea, cosq_val_in_rnea, qd_val_in_rnea, qdd_val_in_rnea,
        v_prev_vec_in_AX_rnea, v_prev_vec_in_AY_rnea, v_prev_vec_in_AZ_rnea, v_prev_vec_in_LX_rnea, v_prev_vec_in_LY_rnea, v_prev_vec_in_LZ_rnea, a_prev_vec_in_AX_rnea, a_prev_vec_in_AY_rnea, a_prev_vec_in_AZ_rnea, a_prev_vec_in_LX_rnea, a_prev_vec_in_LY_rnea, a_prev_vec_in_LZ_rnea,
        link_in_dqPE1, link_in_dqPE2, link_in_dqPE3, link_in_dqPE4, link_in_dqPE5, link_in_dqPE6, link_in_dqPE7, link_in_dqdPE1, link_in_dqdPE2, link_in_dqdPE3, link_in_dqdPE4, link_in_dqdPE5, link_in_dqdPE6, link_in_dqdPE7, derv_in_dqPE1, derv_in_dqPE2, derv_in_dqPE3, derv_in_dqPE4, derv_in_dqPE5, derv_in_dqPE6, derv_in_dqPE7, derv_in_dqdPE1, derv_in_dqdPE2, derv_in_dqdPE3, derv_in_dqdPE4, derv_in_dqdPE5, derv_in_dqdPE6, derv_in_dqdPE7,
        sinq_val_in_dqPE1, sinq_val_in_dqPE2, sinq_val_in_dqPE3, sinq_val_in_dqPE4, sinq_val_in_dqPE5, sinq_val_in_dqPE6, sinq_val_in_dqPE7, sinq_val_in_dqdPE1, sinq_val_in_dqdPE2, sinq_val_in_dqdPE3, sinq_val_in_dqdPE4, sinq_val_in_dqdPE5, sinq_val_in_dqdPE6, sinq_val_in_dqdPE7, cosq_val_in_dqPE1, cosq_val_in_dqPE2, cosq_val_in_dqPE3, cosq_val_in_dqPE4, cosq_val_in_dqPE5, cosq_val_in_dqPE6, cosq_val_in_dqPE7, cosq_val_in_dqdPE1, cosq_val_in_dqdPE2, cosq_val_in_dqdPE3, cosq_val_in_dqdPE4, cosq_val_in_dqdPE5, cosq_val_in_dqdPE6, cosq_val_in_dqdPE7, qd_val_in_dqPE1, qd_val_in_dqPE2, qd_val_in_dqPE3, qd_val_in_dqPE4, qd_val_in_dqPE5, qd_val_in_dqPE6, qd_val_in_dqPE7, qd_val_in_dqdPE1, qd_val_in_dqdPE2, qd_val_in_dqdPE3, qd_val_in_dqdPE4, qd_val_in_dqdPE5, qd_val_in_dqdPE6, qd_val_in_dqdPE7,
        v_curr_vec_in_AX_dqPE1, v_curr_vec_in_AY_dqPE1, v_curr_vec_in_AZ_dqPE1, v_curr_vec_in_LX_dqPE1, v_curr_vec_in_LY_dqPE1, v_curr_vec_in_LZ_dqPE1, v_curr_vec_in_AX_dqPE2, v_curr_vec_in_AY_dqPE2, v_curr_vec_in_AZ_dqPE2, v_curr_vec_in_LX_dqPE2, v_curr_vec_in_LY_dqPE2, v_curr_vec_in_LZ_dqPE2, v_curr_vec_in_AX_dqPE3, v_curr_vec_in_AY_dqPE3, v_curr_vec_in_AZ_dqPE3, v_curr_vec_in_LX_dqPE3, v_curr_vec_in_LY_dqPE3, v_curr_vec_in_LZ_dqPE3, v_curr_vec_in_AX_dqPE4, v_curr_vec_in_AY_dqPE4, v_curr_vec_in_AZ_dqPE4, v_curr_vec_in_LX_dqPE4, v_curr_vec_in_LY_dqPE4, v_curr_vec_in_LZ_dqPE4, v_curr_vec_in_AX_dqPE5, v_curr_vec_in_AY_dqPE5, v_curr_vec_in_AZ_dqPE5, v_curr_vec_in_LX_dqPE5, v_curr_vec_in_LY_dqPE5, v_curr_vec_in_LZ_dqPE5, v_curr_vec_in_AX_dqPE6, v_curr_vec_in_AY_dqPE6, v_curr_vec_in_AZ_dqPE6, v_curr_vec_in_LX_dqPE6, v_curr_vec_in_LY_dqPE6, v_curr_vec_in_LZ_dqPE6, v_curr_vec_in_AX_dqPE7, v_curr_vec_in_AY_dqPE7, v_curr_vec_in_AZ_dqPE7, v_curr_vec_in_LX_dqPE7, v_curr_vec_in_LY_dqPE7, v_curr_vec_in_LZ_dqPE7, v_curr_vec_in_AX_dqdPE1, v_curr_vec_in_AY_dqdPE1, v_curr_vec_in_AZ_dqdPE1, v_curr_vec_in_LX_dqdPE1, v_curr_vec_in_LY_dqdPE1, v_curr_vec_in_LZ_dqdPE1, v_curr_vec_in_AX_dqdPE2, v_curr_vec_in_AY_dqdPE2, v_curr_vec_in_AZ_dqdPE2, v_curr_vec_in_LX_dqdPE2, v_curr_vec_in_LY_dqdPE2, v_curr_vec_in_LZ_dqdPE2, v_curr_vec_in_AX_dqdPE3, v_curr_vec_in_AY_dqdPE3, v_curr_vec_in_AZ_dqdPE3, v_curr_vec_in_LX_dqdPE3, v_curr_vec_in_LY_dqdPE3, v_curr_vec_in_LZ_dqdPE3, v_curr_vec_in_AX_dqdPE4, v_curr_vec_in_AY_dqdPE4, v_curr_vec_in_AZ_dqdPE4, v_curr_vec_in_LX_dqdPE4, v_curr_vec_in_LY_dqdPE4, v_curr_vec_in_LZ_dqdPE4, v_curr_vec_in_AX_dqdPE5, v_curr_vec_in_AY_dqdPE5, v_curr_vec_in_AZ_dqdPE5, v_curr_vec_in_LX_dqdPE5, v_curr_vec_in_LY_dqdPE5, v_curr_vec_in_LZ_dqdPE5, v_curr_vec_in_AX_dqdPE6, v_curr_vec_in_AY_dqdPE6, v_curr_vec_in_AZ_dqdPE6, v_curr_vec_in_LX_dqdPE6, v_curr_vec_in_LY_dqdPE6, v_curr_vec_in_LZ_dqdPE6, v_curr_vec_in_AX_dqdPE7, v_curr_vec_in_AY_dqdPE7, v_curr_vec_in_AZ_dqdPE7, v_curr_vec_in_LX_dqdPE7, v_curr_vec_in_LY_dqdPE7, v_curr_vec_in_LZ_dqdPE7, a_curr_vec_in_AX_dqPE1, a_curr_vec_in_AY_dqPE1, a_curr_vec_in_AZ_dqPE1, a_curr_vec_in_LX_dqPE1, a_curr_vec_in_LY_dqPE1, a_curr_vec_in_LZ_dqPE1, a_curr_vec_in_AX_dqPE2, a_curr_vec_in_AY_dqPE2, a_curr_vec_in_AZ_dqPE2, a_curr_vec_in_LX_dqPE2, a_curr_vec_in_LY_dqPE2, a_curr_vec_in_LZ_dqPE2, a_curr_vec_in_AX_dqPE3, a_curr_vec_in_AY_dqPE3, a_curr_vec_in_AZ_dqPE3, a_curr_vec_in_LX_dqPE3, a_curr_vec_in_LY_dqPE3, a_curr_vec_in_LZ_dqPE3, a_curr_vec_in_AX_dqPE4, a_curr_vec_in_AY_dqPE4, a_curr_vec_in_AZ_dqPE4, a_curr_vec_in_LX_dqPE4, a_curr_vec_in_LY_dqPE4, a_curr_vec_in_LZ_dqPE4, a_curr_vec_in_AX_dqPE5, a_curr_vec_in_AY_dqPE5, a_curr_vec_in_AZ_dqPE5, a_curr_vec_in_LX_dqPE5, a_curr_vec_in_LY_dqPE5, a_curr_vec_in_LZ_dqPE5, a_curr_vec_in_AX_dqPE6, a_curr_vec_in_AY_dqPE6, a_curr_vec_in_AZ_dqPE6, a_curr_vec_in_LX_dqPE6, a_curr_vec_in_LY_dqPE6, a_curr_vec_in_LZ_dqPE6, a_curr_vec_in_AX_dqPE7, a_curr_vec_in_AY_dqPE7, a_curr_vec_in_AZ_dqPE7, a_curr_vec_in_LX_dqPE7, a_curr_vec_in_LY_dqPE7, a_curr_vec_in_LZ_dqPE7, a_curr_vec_in_AX_dqdPE1, a_curr_vec_in_AY_dqdPE1, a_curr_vec_in_AZ_dqdPE1, a_curr_vec_in_LX_dqdPE1, a_curr_vec_in_LY_dqdPE1, a_curr_vec_in_LZ_dqdPE1, a_curr_vec_in_AX_dqdPE2, a_curr_vec_in_AY_dqdPE2, a_curr_vec_in_AZ_dqdPE2, a_curr_vec_in_LX_dqdPE2, a_curr_vec_in_LY_dqdPE2, a_curr_vec_in_LZ_dqdPE2, a_curr_vec_in_AX_dqdPE3, a_curr_vec_in_AY_dqdPE3, a_curr_vec_in_AZ_dqdPE3, a_curr_vec_in_LX_dqdPE3, a_curr_vec_in_LY_dqdPE3, a_curr_vec_in_LZ_dqdPE3, a_curr_vec_in_AX_dqdPE4, a_curr_vec_in_AY_dqdPE4, a_curr_vec_in_AZ_dqdPE4, a_curr_vec_in_LX_dqdPE4, a_curr_vec_in_LY_dqdPE4, a_curr_vec_in_LZ_dqdPE4, a_curr_vec_in_AX_dqdPE5, a_curr_vec_in_AY_dqdPE5, a_curr_vec_in_AZ_dqdPE5, a_curr_vec_in_LX_dqdPE5, a_curr_vec_in_LY_dqdPE5, a_curr_vec_in_LZ_dqdPE5, a_curr_vec_in_AX_dqdPE6, a_curr_vec_in_AY_dqdPE6, a_curr_vec_in_AZ_dqdPE6, a_curr_vec_in_LX_dqdPE6, a_curr_vec_in_LY_dqdPE6, a_curr_vec_in_LZ_dqdPE6, a_curr_vec_in_AX_dqdPE7, a_curr_vec_in_AY_dqdPE7, a_curr_vec_in_AZ_dqdPE7, a_curr_vec_in_LX_dqdPE7, a_curr_vec_in_LY_dqdPE7, a_curr_vec_in_LZ_dqdPE7, v_prev_vec_in_AX_dqPE1, v_prev_vec_in_AY_dqPE1, v_prev_vec_in_AZ_dqPE1, v_prev_vec_in_LX_dqPE1, v_prev_vec_in_LY_dqPE1, v_prev_vec_in_LZ_dqPE1, v_prev_vec_in_AX_dqPE2, v_prev_vec_in_AY_dqPE2, v_prev_vec_in_AZ_dqPE2, v_prev_vec_in_LX_dqPE2, v_prev_vec_in_LY_dqPE2, v_prev_vec_in_LZ_dqPE2, v_prev_vec_in_AX_dqPE3, v_prev_vec_in_AY_dqPE3, v_prev_vec_in_AZ_dqPE3, v_prev_vec_in_LX_dqPE3, v_prev_vec_in_LY_dqPE3, v_prev_vec_in_LZ_dqPE3, v_prev_vec_in_AX_dqPE4, v_prev_vec_in_AY_dqPE4, v_prev_vec_in_AZ_dqPE4, v_prev_vec_in_LX_dqPE4, v_prev_vec_in_LY_dqPE4, v_prev_vec_in_LZ_dqPE4, v_prev_vec_in_AX_dqPE5, v_prev_vec_in_AY_dqPE5, v_prev_vec_in_AZ_dqPE5, v_prev_vec_in_LX_dqPE5, v_prev_vec_in_LY_dqPE5, v_prev_vec_in_LZ_dqPE5, v_prev_vec_in_AX_dqPE6, v_prev_vec_in_AY_dqPE6, v_prev_vec_in_AZ_dqPE6, v_prev_vec_in_LX_dqPE6, v_prev_vec_in_LY_dqPE6, v_prev_vec_in_LZ_dqPE6, v_prev_vec_in_AX_dqPE7, v_prev_vec_in_AY_dqPE7, v_prev_vec_in_AZ_dqPE7, v_prev_vec_in_LX_dqPE7, v_prev_vec_in_LY_dqPE7, v_prev_vec_in_LZ_dqPE7, a_prev_vec_in_AX_dqPE1, a_prev_vec_in_AY_dqPE1, a_prev_vec_in_AZ_dqPE1, a_prev_vec_in_LX_dqPE1, a_prev_vec_in_LY_dqPE1, a_prev_vec_in_LZ_dqPE1, a_prev_vec_in_AX_dqPE2, a_prev_vec_in_AY_dqPE2, a_prev_vec_in_AZ_dqPE2, a_prev_vec_in_LX_dqPE2, a_prev_vec_in_LY_dqPE2, a_prev_vec_in_LZ_dqPE2, a_prev_vec_in_AX_dqPE3, a_prev_vec_in_AY_dqPE3, a_prev_vec_in_AZ_dqPE3, a_prev_vec_in_LX_dqPE3, a_prev_vec_in_LY_dqPE3, a_prev_vec_in_LZ_dqPE3, a_prev_vec_in_AX_dqPE4, a_prev_vec_in_AY_dqPE4, a_prev_vec_in_AZ_dqPE4, a_prev_vec_in_LX_dqPE4, a_prev_vec_in_LY_dqPE4, a_prev_vec_in_LZ_dqPE4, a_prev_vec_in_AX_dqPE5, a_prev_vec_in_AY_dqPE5, a_prev_vec_in_AZ_dqPE5, a_prev_vec_in_LX_dqPE5, a_prev_vec_in_LY_dqPE5, a_prev_vec_in_LZ_dqPE5, a_prev_vec_in_AX_dqPE6, a_prev_vec_in_AY_dqPE6, a_prev_vec_in_AZ_dqPE6, a_prev_vec_in_LX_dqPE6, a_prev_vec_in_LY_dqPE6, a_prev_vec_in_LZ_dqPE6, a_prev_vec_in_AX_dqPE7, a_prev_vec_in_AY_dqPE7, a_prev_vec_in_AZ_dqPE7, a_prev_vec_in_LX_dqPE7, a_prev_vec_in_LY_dqPE7, a_prev_vec_in_LZ_dqPE7,
        dvdq_prev_vec_in_AX_dqPE1, dvdq_prev_vec_in_AY_dqPE1, dvdq_prev_vec_in_AZ_dqPE1, dvdq_prev_vec_in_LX_dqPE1, dvdq_prev_vec_in_LY_dqPE1, dvdq_prev_vec_in_LZ_dqPE1, dvdq_prev_vec_in_AX_dqPE2, dvdq_prev_vec_in_AY_dqPE2, dvdq_prev_vec_in_AZ_dqPE2, dvdq_prev_vec_in_LX_dqPE2, dvdq_prev_vec_in_LY_dqPE2, dvdq_prev_vec_in_LZ_dqPE2, dvdq_prev_vec_in_AX_dqPE3, dvdq_prev_vec_in_AY_dqPE3, dvdq_prev_vec_in_AZ_dqPE3, dvdq_prev_vec_in_LX_dqPE3, dvdq_prev_vec_in_LY_dqPE3, dvdq_prev_vec_in_LZ_dqPE3, dvdq_prev_vec_in_AX_dqPE4, dvdq_prev_vec_in_AY_dqPE4, dvdq_prev_vec_in_AZ_dqPE4, dvdq_prev_vec_in_LX_dqPE4, dvdq_prev_vec_in_LY_dqPE4, dvdq_prev_vec_in_LZ_dqPE4, dvdq_prev_vec_in_AX_dqPE5, dvdq_prev_vec_in_AY_dqPE5, dvdq_prev_vec_in_AZ_dqPE5, dvdq_prev_vec_in_LX_dqPE5, dvdq_prev_vec_in_LY_dqPE5, dvdq_prev_vec_in_LZ_dqPE5, dvdq_prev_vec_in_AX_dqPE6, dvdq_prev_vec_in_AY_dqPE6, dvdq_prev_vec_in_AZ_dqPE6, dvdq_prev_vec_in_LX_dqPE6, dvdq_prev_vec_in_LY_dqPE6, dvdq_prev_vec_in_LZ_dqPE6, dvdq_prev_vec_in_AX_dqPE7, dvdq_prev_vec_in_AY_dqPE7, dvdq_prev_vec_in_AZ_dqPE7, dvdq_prev_vec_in_LX_dqPE7, dvdq_prev_vec_in_LY_dqPE7, dvdq_prev_vec_in_LZ_dqPE7, dvdqd_prev_vec_in_AX_dqdPE1, dvdqd_prev_vec_in_AY_dqdPE1, dvdqd_prev_vec_in_AZ_dqdPE1, dvdqd_prev_vec_in_LX_dqdPE1, dvdqd_prev_vec_in_LY_dqdPE1, dvdqd_prev_vec_in_LZ_dqdPE1, dvdqd_prev_vec_in_AX_dqdPE2, dvdqd_prev_vec_in_AY_dqdPE2, dvdqd_prev_vec_in_AZ_dqdPE2, dvdqd_prev_vec_in_LX_dqdPE2, dvdqd_prev_vec_in_LY_dqdPE2, dvdqd_prev_vec_in_LZ_dqdPE2, dvdqd_prev_vec_in_AX_dqdPE3, dvdqd_prev_vec_in_AY_dqdPE3, dvdqd_prev_vec_in_AZ_dqdPE3, dvdqd_prev_vec_in_LX_dqdPE3, dvdqd_prev_vec_in_LY_dqdPE3, dvdqd_prev_vec_in_LZ_dqdPE3, dvdqd_prev_vec_in_AX_dqdPE4, dvdqd_prev_vec_in_AY_dqdPE4, dvdqd_prev_vec_in_AZ_dqdPE4, dvdqd_prev_vec_in_LX_dqdPE4, dvdqd_prev_vec_in_LY_dqdPE4, dvdqd_prev_vec_in_LZ_dqdPE4, dvdqd_prev_vec_in_AX_dqdPE5, dvdqd_prev_vec_in_AY_dqdPE5, dvdqd_prev_vec_in_AZ_dqdPE5, dvdqd_prev_vec_in_LX_dqdPE5, dvdqd_prev_vec_in_LY_dqdPE5, dvdqd_prev_vec_in_LZ_dqdPE5, dvdqd_prev_vec_in_AX_dqdPE6, dvdqd_prev_vec_in_AY_dqdPE6, dvdqd_prev_vec_in_AZ_dqdPE6, dvdqd_prev_vec_in_LX_dqdPE6, dvdqd_prev_vec_in_LY_dqdPE6, dvdqd_prev_vec_in_LZ_dqdPE6, dvdqd_prev_vec_in_AX_dqdPE7, dvdqd_prev_vec_in_AY_dqdPE7, dvdqd_prev_vec_in_AZ_dqdPE7, dvdqd_prev_vec_in_LX_dqdPE7, dvdqd_prev_vec_in_LY_dqdPE7, dvdqd_prev_vec_in_LZ_dqdPE7, dadq_prev_vec_in_AX_dqPE1, dadq_prev_vec_in_AY_dqPE1, dadq_prev_vec_in_AZ_dqPE1, dadq_prev_vec_in_LX_dqPE1, dadq_prev_vec_in_LY_dqPE1, dadq_prev_vec_in_LZ_dqPE1, dadq_prev_vec_in_AX_dqPE2, dadq_prev_vec_in_AY_dqPE2, dadq_prev_vec_in_AZ_dqPE2, dadq_prev_vec_in_LX_dqPE2, dadq_prev_vec_in_LY_dqPE2, dadq_prev_vec_in_LZ_dqPE2, dadq_prev_vec_in_AX_dqPE3, dadq_prev_vec_in_AY_dqPE3, dadq_prev_vec_in_AZ_dqPE3, dadq_prev_vec_in_LX_dqPE3, dadq_prev_vec_in_LY_dqPE3, dadq_prev_vec_in_LZ_dqPE3, dadq_prev_vec_in_AX_dqPE4, dadq_prev_vec_in_AY_dqPE4, dadq_prev_vec_in_AZ_dqPE4, dadq_prev_vec_in_LX_dqPE4, dadq_prev_vec_in_LY_dqPE4, dadq_prev_vec_in_LZ_dqPE4, dadq_prev_vec_in_AX_dqPE5, dadq_prev_vec_in_AY_dqPE5, dadq_prev_vec_in_AZ_dqPE5, dadq_prev_vec_in_LX_dqPE5, dadq_prev_vec_in_LY_dqPE5, dadq_prev_vec_in_LZ_dqPE5, dadq_prev_vec_in_AX_dqPE6, dadq_prev_vec_in_AY_dqPE6, dadq_prev_vec_in_AZ_dqPE6, dadq_prev_vec_in_LX_dqPE6, dadq_prev_vec_in_LY_dqPE6, dadq_prev_vec_in_LZ_dqPE6, dadq_prev_vec_in_AX_dqPE7, dadq_prev_vec_in_AY_dqPE7, dadq_prev_vec_in_AZ_dqPE7, dadq_prev_vec_in_LX_dqPE7, dadq_prev_vec_in_LY_dqPE7, dadq_prev_vec_in_LZ_dqPE7, dadqd_prev_vec_in_AX_dqdPE1, dadqd_prev_vec_in_AY_dqdPE1, dadqd_prev_vec_in_AZ_dqdPE1, dadqd_prev_vec_in_LX_dqdPE1, dadqd_prev_vec_in_LY_dqdPE1, dadqd_prev_vec_in_LZ_dqdPE1, dadqd_prev_vec_in_AX_dqdPE2, dadqd_prev_vec_in_AY_dqdPE2, dadqd_prev_vec_in_AZ_dqdPE2, dadqd_prev_vec_in_LX_dqdPE2, dadqd_prev_vec_in_LY_dqdPE2, dadqd_prev_vec_in_LZ_dqdPE2, dadqd_prev_vec_in_AX_dqdPE3, dadqd_prev_vec_in_AY_dqdPE3, dadqd_prev_vec_in_AZ_dqdPE3, dadqd_prev_vec_in_LX_dqdPE3, dadqd_prev_vec_in_LY_dqdPE3, dadqd_prev_vec_in_LZ_dqdPE3, dadqd_prev_vec_in_AX_dqdPE4, dadqd_prev_vec_in_AY_dqdPE4, dadqd_prev_vec_in_AZ_dqdPE4, dadqd_prev_vec_in_LX_dqdPE4, dadqd_prev_vec_in_LY_dqdPE4, dadqd_prev_vec_in_LZ_dqdPE4, dadqd_prev_vec_in_AX_dqdPE5, dadqd_prev_vec_in_AY_dqdPE5, dadqd_prev_vec_in_AZ_dqdPE5, dadqd_prev_vec_in_LX_dqdPE5, dadqd_prev_vec_in_LY_dqdPE5, dadqd_prev_vec_in_LZ_dqdPE5, dadqd_prev_vec_in_AX_dqdPE6, dadqd_prev_vec_in_AY_dqdPE6, dadqd_prev_vec_in_AZ_dqdPE6, dadqd_prev_vec_in_LX_dqdPE6, dadqd_prev_vec_in_LY_dqdPE6, dadqd_prev_vec_in_LZ_dqdPE6, dadqd_prev_vec_in_AX_dqdPE7, dadqd_prev_vec_in_AY_dqdPE7, dadqd_prev_vec_in_AZ_dqdPE7, dadqd_prev_vec_in_LX_dqdPE7, dadqd_prev_vec_in_LY_dqdPE7, dadqd_prev_vec_in_LZ_dqdPE7,
        output_ready,
        v_curr_vec_out_AX_rnea, v_curr_vec_out_AY_rnea, v_curr_vec_out_AZ_rnea, v_curr_vec_out_LX_rnea, v_curr_vec_out_LY_rnea, v_curr_vec_out_LZ_rnea, a_curr_vec_out_AX_rnea, a_curr_vec_out_AY_rnea, a_curr_vec_out_AZ_rnea, a_curr_vec_out_LX_rnea, a_curr_vec_out_LY_rnea, a_curr_vec_out_LZ_rnea, f_curr_vec_out_AX_rnea, f_curr_vec_out_AY_rnea, f_curr_vec_out_AZ_rnea, f_curr_vec_out_LX_rnea, f_curr_vec_out_LY_rnea, f_curr_vec_out_LZ_rnea,
        dfdq_curr_vec_out_AX_dqPE1, dfdq_curr_vec_out_AY_dqPE1, dfdq_curr_vec_out_AZ_dqPE1, dfdq_curr_vec_out_LX_dqPE1, dfdq_curr_vec_out_LY_dqPE1, dfdq_curr_vec_out_LZ_dqPE1, dfdq_curr_vec_out_AX_dqPE2, dfdq_curr_vec_out_AY_dqPE2, dfdq_curr_vec_out_AZ_dqPE2, dfdq_curr_vec_out_LX_dqPE2, dfdq_curr_vec_out_LY_dqPE2, dfdq_curr_vec_out_LZ_dqPE2, dfdq_curr_vec_out_AX_dqPE3, dfdq_curr_vec_out_AY_dqPE3, dfdq_curr_vec_out_AZ_dqPE3, dfdq_curr_vec_out_LX_dqPE3, dfdq_curr_vec_out_LY_dqPE3, dfdq_curr_vec_out_LZ_dqPE3, dfdq_curr_vec_out_AX_dqPE4, dfdq_curr_vec_out_AY_dqPE4, dfdq_curr_vec_out_AZ_dqPE4, dfdq_curr_vec_out_LX_dqPE4, dfdq_curr_vec_out_LY_dqPE4, dfdq_curr_vec_out_LZ_dqPE4, dfdq_curr_vec_out_AX_dqPE5, dfdq_curr_vec_out_AY_dqPE5, dfdq_curr_vec_out_AZ_dqPE5, dfdq_curr_vec_out_LX_dqPE5, dfdq_curr_vec_out_LY_dqPE5, dfdq_curr_vec_out_LZ_dqPE5, dfdq_curr_vec_out_AX_dqPE6, dfdq_curr_vec_out_AY_dqPE6, dfdq_curr_vec_out_AZ_dqPE6, dfdq_curr_vec_out_LX_dqPE6, dfdq_curr_vec_out_LY_dqPE6, dfdq_curr_vec_out_LZ_dqPE6, dfdq_curr_vec_out_AX_dqPE7, dfdq_curr_vec_out_AY_dqPE7, dfdq_curr_vec_out_AZ_dqPE7, dfdq_curr_vec_out_LX_dqPE7, dfdq_curr_vec_out_LY_dqPE7, dfdq_curr_vec_out_LZ_dqPE7, dfdqd_curr_vec_out_AX_dqdPE1, dfdqd_curr_vec_out_AY_dqdPE1, dfdqd_curr_vec_out_AZ_dqdPE1, dfdqd_curr_vec_out_LX_dqdPE1, dfdqd_curr_vec_out_LY_dqdPE1, dfdqd_curr_vec_out_LZ_dqdPE1, dfdqd_curr_vec_out_AX_dqdPE2, dfdqd_curr_vec_out_AY_dqdPE2, dfdqd_curr_vec_out_AZ_dqdPE2, dfdqd_curr_vec_out_LX_dqdPE2, dfdqd_curr_vec_out_LY_dqdPE2, dfdqd_curr_vec_out_LZ_dqdPE2, dfdqd_curr_vec_out_AX_dqdPE3, dfdqd_curr_vec_out_AY_dqdPE3, dfdqd_curr_vec_out_AZ_dqdPE3, dfdqd_curr_vec_out_LX_dqdPE3, dfdqd_curr_vec_out_LY_dqdPE3, dfdqd_curr_vec_out_LZ_dqdPE3, dfdqd_curr_vec_out_AX_dqdPE4, dfdqd_curr_vec_out_AY_dqdPE4, dfdqd_curr_vec_out_AZ_dqdPE4, dfdqd_curr_vec_out_LX_dqdPE4, dfdqd_curr_vec_out_LY_dqdPE4, dfdqd_curr_vec_out_LZ_dqdPE4, dfdqd_curr_vec_out_AX_dqdPE5, dfdqd_curr_vec_out_AY_dqdPE5, dfdqd_curr_vec_out_AZ_dqdPE5, dfdqd_curr_vec_out_LX_dqdPE5, dfdqd_curr_vec_out_LY_dqdPE5, dfdqd_curr_vec_out_LZ_dqdPE5, dfdqd_curr_vec_out_AX_dqdPE6, dfdqd_curr_vec_out_AY_dqdPE6, dfdqd_curr_vec_out_AZ_dqdPE6, dfdqd_curr_vec_out_LX_dqdPE6, dfdqd_curr_vec_out_LY_dqdPE6, dfdqd_curr_vec_out_LZ_dqdPE6, dfdqd_curr_vec_out_AX_dqdPE7, dfdqd_curr_vec_out_AY_dqdPE7, dfdqd_curr_vec_out_AZ_dqdPE7, dfdqd_curr_vec_out_LX_dqdPE7, dfdqd_curr_vec_out_LY_dqdPE7, dfdqd_curr_vec_out_LZ_dqdPE7,
        dvdq_curr_vec_out_AX_dqPE1, dvdq_curr_vec_out_AY_dqPE1, dvdq_curr_vec_out_AZ_dqPE1, dvdq_curr_vec_out_LX_dqPE1, dvdq_curr_vec_out_LY_dqPE1, dvdq_curr_vec_out_LZ_dqPE1, dvdq_curr_vec_out_AX_dqPE2, dvdq_curr_vec_out_AY_dqPE2, dvdq_curr_vec_out_AZ_dqPE2, dvdq_curr_vec_out_LX_dqPE2, dvdq_curr_vec_out_LY_dqPE2, dvdq_curr_vec_out_LZ_dqPE2, dvdq_curr_vec_out_AX_dqPE3, dvdq_curr_vec_out_AY_dqPE3, dvdq_curr_vec_out_AZ_dqPE3, dvdq_curr_vec_out_LX_dqPE3, dvdq_curr_vec_out_LY_dqPE3, dvdq_curr_vec_out_LZ_dqPE3, dvdq_curr_vec_out_AX_dqPE4, dvdq_curr_vec_out_AY_dqPE4, dvdq_curr_vec_out_AZ_dqPE4, dvdq_curr_vec_out_LX_dqPE4, dvdq_curr_vec_out_LY_dqPE4, dvdq_curr_vec_out_LZ_dqPE4, dvdq_curr_vec_out_AX_dqPE5, dvdq_curr_vec_out_AY_dqPE5, dvdq_curr_vec_out_AZ_dqPE5, dvdq_curr_vec_out_LX_dqPE5, dvdq_curr_vec_out_LY_dqPE5, dvdq_curr_vec_out_LZ_dqPE5, dvdq_curr_vec_out_AX_dqPE6, dvdq_curr_vec_out_AY_dqPE6, dvdq_curr_vec_out_AZ_dqPE6, dvdq_curr_vec_out_LX_dqPE6, dvdq_curr_vec_out_LY_dqPE6, dvdq_curr_vec_out_LZ_dqPE6, dvdq_curr_vec_out_AX_dqPE7, dvdq_curr_vec_out_AY_dqPE7, dvdq_curr_vec_out_AZ_dqPE7, dvdq_curr_vec_out_LX_dqPE7, dvdq_curr_vec_out_LY_dqPE7, dvdq_curr_vec_out_LZ_dqPE7, dvdqd_curr_vec_out_AX_dqdPE1, dvdqd_curr_vec_out_AY_dqdPE1, dvdqd_curr_vec_out_AZ_dqdPE1, dvdqd_curr_vec_out_LX_dqdPE1, dvdqd_curr_vec_out_LY_dqdPE1, dvdqd_curr_vec_out_LZ_dqdPE1, dvdqd_curr_vec_out_AX_dqdPE2, dvdqd_curr_vec_out_AY_dqdPE2, dvdqd_curr_vec_out_AZ_dqdPE2, dvdqd_curr_vec_out_LX_dqdPE2, dvdqd_curr_vec_out_LY_dqdPE2, dvdqd_curr_vec_out_LZ_dqdPE2, dvdqd_curr_vec_out_AX_dqdPE3, dvdqd_curr_vec_out_AY_dqdPE3, dvdqd_curr_vec_out_AZ_dqdPE3, dvdqd_curr_vec_out_LX_dqdPE3, dvdqd_curr_vec_out_LY_dqdPE3, dvdqd_curr_vec_out_LZ_dqdPE3, dvdqd_curr_vec_out_AX_dqdPE4, dvdqd_curr_vec_out_AY_dqdPE4, dvdqd_curr_vec_out_AZ_dqdPE4, dvdqd_curr_vec_out_LX_dqdPE4, dvdqd_curr_vec_out_LY_dqdPE4, dvdqd_curr_vec_out_LZ_dqdPE4, dvdqd_curr_vec_out_AX_dqdPE5, dvdqd_curr_vec_out_AY_dqdPE5, dvdqd_curr_vec_out_AZ_dqdPE5, dvdqd_curr_vec_out_LX_dqdPE5, dvdqd_curr_vec_out_LY_dqdPE5, dvdqd_curr_vec_out_LZ_dqdPE5, dvdqd_curr_vec_out_AX_dqdPE6, dvdqd_curr_vec_out_AY_dqdPE6, dvdqd_curr_vec_out_AZ_dqdPE6, dvdqd_curr_vec_out_LX_dqdPE6, dvdqd_curr_vec_out_LY_dqdPE6, dvdqd_curr_vec_out_LZ_dqdPE6, dvdqd_curr_vec_out_AX_dqdPE7, dvdqd_curr_vec_out_AY_dqdPE7, dvdqd_curr_vec_out_AZ_dqdPE7, dvdqd_curr_vec_out_LX_dqdPE7, dvdqd_curr_vec_out_LY_dqdPE7, dvdqd_curr_vec_out_LZ_dqdPE7, dadq_curr_vec_out_AX_dqPE1, dadq_curr_vec_out_AY_dqPE1, dadq_curr_vec_out_AZ_dqPE1, dadq_curr_vec_out_LX_dqPE1, dadq_curr_vec_out_LY_dqPE1, dadq_curr_vec_out_LZ_dqPE1, dadq_curr_vec_out_AX_dqPE2, dadq_curr_vec_out_AY_dqPE2, dadq_curr_vec_out_AZ_dqPE2, dadq_curr_vec_out_LX_dqPE2, dadq_curr_vec_out_LY_dqPE2, dadq_curr_vec_out_LZ_dqPE2, dadq_curr_vec_out_AX_dqPE3, dadq_curr_vec_out_AY_dqPE3, dadq_curr_vec_out_AZ_dqPE3, dadq_curr_vec_out_LX_dqPE3, dadq_curr_vec_out_LY_dqPE3, dadq_curr_vec_out_LZ_dqPE3, dadq_curr_vec_out_AX_dqPE4, dadq_curr_vec_out_AY_dqPE4, dadq_curr_vec_out_AZ_dqPE4, dadq_curr_vec_out_LX_dqPE4, dadq_curr_vec_out_LY_dqPE4, dadq_curr_vec_out_LZ_dqPE4, dadq_curr_vec_out_AX_dqPE5, dadq_curr_vec_out_AY_dqPE5, dadq_curr_vec_out_AZ_dqPE5, dadq_curr_vec_out_LX_dqPE5, dadq_curr_vec_out_LY_dqPE5, dadq_curr_vec_out_LZ_dqPE5, dadq_curr_vec_out_AX_dqPE6, dadq_curr_vec_out_AY_dqPE6, dadq_curr_vec_out_AZ_dqPE6, dadq_curr_vec_out_LX_dqPE6, dadq_curr_vec_out_LY_dqPE6, dadq_curr_vec_out_LZ_dqPE6, dadq_curr_vec_out_AX_dqPE7, dadq_curr_vec_out_AY_dqPE7, dadq_curr_vec_out_AZ_dqPE7, dadq_curr_vec_out_LX_dqPE7, dadq_curr_vec_out_LY_dqPE7, dadq_curr_vec_out_LZ_dqPE7, dadqd_curr_vec_out_AX_dqdPE1, dadqd_curr_vec_out_AY_dqdPE1, dadqd_curr_vec_out_AZ_dqdPE1, dadqd_curr_vec_out_LX_dqdPE1, dadqd_curr_vec_out_LY_dqdPE1, dadqd_curr_vec_out_LZ_dqdPE1, dadqd_curr_vec_out_AX_dqdPE2, dadqd_curr_vec_out_AY_dqdPE2, dadqd_curr_vec_out_AZ_dqdPE2, dadqd_curr_vec_out_LX_dqdPE2, dadqd_curr_vec_out_LY_dqdPE2, dadqd_curr_vec_out_LZ_dqdPE2, dadqd_curr_vec_out_AX_dqdPE3, dadqd_curr_vec_out_AY_dqdPE3, dadqd_curr_vec_out_AZ_dqdPE3, dadqd_curr_vec_out_LX_dqdPE3, dadqd_curr_vec_out_LY_dqdPE3, dadqd_curr_vec_out_LZ_dqdPE3, dadqd_curr_vec_out_AX_dqdPE4, dadqd_curr_vec_out_AY_dqdPE4, dadqd_curr_vec_out_AZ_dqdPE4, dadqd_curr_vec_out_LX_dqdPE4, dadqd_curr_vec_out_LY_dqdPE4, dadqd_curr_vec_out_LZ_dqdPE4, dadqd_curr_vec_out_AX_dqdPE5, dadqd_curr_vec_out_AY_dqdPE5, dadqd_curr_vec_out_AZ_dqdPE5, dadqd_curr_vec_out_LX_dqdPE5, dadqd_curr_vec_out_LY_dqdPE5, dadqd_curr_vec_out_LZ_dqdPE5, dadqd_curr_vec_out_AX_dqdPE6, dadqd_curr_vec_out_AY_dqdPE6, dadqd_curr_vec_out_AZ_dqdPE6, dadqd_curr_vec_out_LX_dqdPE6, dadqd_curr_vec_out_LY_dqdPE6, dadqd_curr_vec_out_LZ_dqdPE6, dadqd_curr_vec_out_AX_dqdPE7, dadqd_curr_vec_out_AY_dqdPE7, dadqd_curr_vec_out_AZ_dqdPE7, dadqd_curr_vec_out_LX_dqdPE7, dadqd_curr_vec_out_LY_dqdPE7, dadqd_curr_vec_out_LZ_dqdPE7
    ) CF (
        get_data, link_in_rnea, sinq_val_in_rnea, cosq_val_in_rnea, qd_val_in_rnea, qdd_val_in_rnea,
        v_prev_vec_in_AX_rnea, v_prev_vec_in_AY_rnea, v_prev_vec_in_AZ_rnea, v_prev_vec_in_LX_rnea, v_prev_vec_in_LY_rnea, v_prev_vec_in_LZ_rnea, a_prev_vec_in_AX_rnea, a_prev_vec_in_AY_rnea, a_prev_vec_in_AZ_rnea, a_prev_vec_in_LX_rnea, a_prev_vec_in_LY_rnea, a_prev_vec_in_LZ_rnea,
        link_in_dqPE1, link_in_dqPE2, link_in_dqPE3, link_in_dqPE4, link_in_dqPE5, link_in_dqPE6, link_in_dqPE7, link_in_dqdPE1, link_in_dqdPE2, link_in_dqdPE3, link_in_dqdPE4, link_in_dqdPE5, link_in_dqdPE6, link_in_dqdPE7, derv_in_dqPE1, derv_in_dqPE2, derv_in_dqPE3, derv_in_dqPE4, derv_in_dqPE5, derv_in_dqPE6, derv_in_dqPE7, derv_in_dqdPE1, derv_in_dqdPE2, derv_in_dqdPE3, derv_in_dqdPE4, derv_in_dqdPE5, derv_in_dqdPE6, derv_in_dqdPE7,
        sinq_val_in_dqPE1, sinq_val_in_dqPE2, sinq_val_in_dqPE3, sinq_val_in_dqPE4, sinq_val_in_dqPE5, sinq_val_in_dqPE6, sinq_val_in_dqPE7, sinq_val_in_dqdPE1, sinq_val_in_dqdPE2, sinq_val_in_dqdPE3, sinq_val_in_dqdPE4, sinq_val_in_dqdPE5, sinq_val_in_dqdPE6, sinq_val_in_dqdPE7, cosq_val_in_dqPE1, cosq_val_in_dqPE2, cosq_val_in_dqPE3, cosq_val_in_dqPE4, cosq_val_in_dqPE5, cosq_val_in_dqPE6, cosq_val_in_dqPE7, cosq_val_in_dqdPE1, cosq_val_in_dqdPE2, cosq_val_in_dqdPE3, cosq_val_in_dqdPE4, cosq_val_in_dqdPE5, cosq_val_in_dqdPE6, cosq_val_in_dqdPE7, qd_val_in_dqPE1, qd_val_in_dqPE2, qd_val_in_dqPE3, qd_val_in_dqPE4, qd_val_in_dqPE5, qd_val_in_dqPE6, qd_val_in_dqPE7, qd_val_in_dqdPE1, qd_val_in_dqdPE2, qd_val_in_dqdPE3, qd_val_in_dqdPE4, qd_val_in_dqdPE5, qd_val_in_dqdPE6, qd_val_in_dqdPE7,
        v_curr_vec_in_AX_dqPE1, v_curr_vec_in_AY_dqPE1, v_curr_vec_in_AZ_dqPE1, v_curr_vec_in_LX_dqPE1, v_curr_vec_in_LY_dqPE1, v_curr_vec_in_LZ_dqPE1, v_curr_vec_in_AX_dqPE2, v_curr_vec_in_AY_dqPE2, v_curr_vec_in_AZ_dqPE2, v_curr_vec_in_LX_dqPE2, v_curr_vec_in_LY_dqPE2, v_curr_vec_in_LZ_dqPE2, v_curr_vec_in_AX_dqPE3, v_curr_vec_in_AY_dqPE3, v_curr_vec_in_AZ_dqPE3, v_curr_vec_in_LX_dqPE3, v_curr_vec_in_LY_dqPE3, v_curr_vec_in_LZ_dqPE3, v_curr_vec_in_AX_dqPE4, v_curr_vec_in_AY_dqPE4, v_curr_vec_in_AZ_dqPE4, v_curr_vec_in_LX_dqPE4, v_curr_vec_in_LY_dqPE4, v_curr_vec_in_LZ_dqPE4, v_curr_vec_in_AX_dqPE5, v_curr_vec_in_AY_dqPE5, v_curr_vec_in_AZ_dqPE5, v_curr_vec_in_LX_dqPE5, v_curr_vec_in_LY_dqPE5, v_curr_vec_in_LZ_dqPE5, v_curr_vec_in_AX_dqPE6, v_curr_vec_in_AY_dqPE6, v_curr_vec_in_AZ_dqPE6, v_curr_vec_in_LX_dqPE6, v_curr_vec_in_LY_dqPE6, v_curr_vec_in_LZ_dqPE6, v_curr_vec_in_AX_dqPE7, v_curr_vec_in_AY_dqPE7, v_curr_vec_in_AZ_dqPE7, v_curr_vec_in_LX_dqPE7, v_curr_vec_in_LY_dqPE7, v_curr_vec_in_LZ_dqPE7, v_curr_vec_in_AX_dqdPE1, v_curr_vec_in_AY_dqdPE1, v_curr_vec_in_AZ_dqdPE1, v_curr_vec_in_LX_dqdPE1, v_curr_vec_in_LY_dqdPE1, v_curr_vec_in_LZ_dqdPE1, v_curr_vec_in_AX_dqdPE2, v_curr_vec_in_AY_dqdPE2, v_curr_vec_in_AZ_dqdPE2, v_curr_vec_in_LX_dqdPE2, v_curr_vec_in_LY_dqdPE2, v_curr_vec_in_LZ_dqdPE2, v_curr_vec_in_AX_dqdPE3, v_curr_vec_in_AY_dqdPE3, v_curr_vec_in_AZ_dqdPE3, v_curr_vec_in_LX_dqdPE3, v_curr_vec_in_LY_dqdPE3, v_curr_vec_in_LZ_dqdPE3, v_curr_vec_in_AX_dqdPE4, v_curr_vec_in_AY_dqdPE4, v_curr_vec_in_AZ_dqdPE4, v_curr_vec_in_LX_dqdPE4, v_curr_vec_in_LY_dqdPE4, v_curr_vec_in_LZ_dqdPE4, v_curr_vec_in_AX_dqdPE5, v_curr_vec_in_AY_dqdPE5, v_curr_vec_in_AZ_dqdPE5, v_curr_vec_in_LX_dqdPE5, v_curr_vec_in_LY_dqdPE5, v_curr_vec_in_LZ_dqdPE5, v_curr_vec_in_AX_dqdPE6, v_curr_vec_in_AY_dqdPE6, v_curr_vec_in_AZ_dqdPE6, v_curr_vec_in_LX_dqdPE6, v_curr_vec_in_LY_dqdPE6, v_curr_vec_in_LZ_dqdPE6, v_curr_vec_in_AX_dqdPE7, v_curr_vec_in_AY_dqdPE7, v_curr_vec_in_AZ_dqdPE7, v_curr_vec_in_LX_dqdPE7, v_curr_vec_in_LY_dqdPE7, v_curr_vec_in_LZ_dqdPE7, a_curr_vec_in_AX_dqPE1, a_curr_vec_in_AY_dqPE1, a_curr_vec_in_AZ_dqPE1, a_curr_vec_in_LX_dqPE1, a_curr_vec_in_LY_dqPE1, a_curr_vec_in_LZ_dqPE1, a_curr_vec_in_AX_dqPE2, a_curr_vec_in_AY_dqPE2, a_curr_vec_in_AZ_dqPE2, a_curr_vec_in_LX_dqPE2, a_curr_vec_in_LY_dqPE2, a_curr_vec_in_LZ_dqPE2, a_curr_vec_in_AX_dqPE3, a_curr_vec_in_AY_dqPE3, a_curr_vec_in_AZ_dqPE3, a_curr_vec_in_LX_dqPE3, a_curr_vec_in_LY_dqPE3, a_curr_vec_in_LZ_dqPE3, a_curr_vec_in_AX_dqPE4, a_curr_vec_in_AY_dqPE4, a_curr_vec_in_AZ_dqPE4, a_curr_vec_in_LX_dqPE4, a_curr_vec_in_LY_dqPE4, a_curr_vec_in_LZ_dqPE4, a_curr_vec_in_AX_dqPE5, a_curr_vec_in_AY_dqPE5, a_curr_vec_in_AZ_dqPE5, a_curr_vec_in_LX_dqPE5, a_curr_vec_in_LY_dqPE5, a_curr_vec_in_LZ_dqPE5, a_curr_vec_in_AX_dqPE6, a_curr_vec_in_AY_dqPE6, a_curr_vec_in_AZ_dqPE6, a_curr_vec_in_LX_dqPE6, a_curr_vec_in_LY_dqPE6, a_curr_vec_in_LZ_dqPE6, a_curr_vec_in_AX_dqPE7, a_curr_vec_in_AY_dqPE7, a_curr_vec_in_AZ_dqPE7, a_curr_vec_in_LX_dqPE7, a_curr_vec_in_LY_dqPE7, a_curr_vec_in_LZ_dqPE7, a_curr_vec_in_AX_dqdPE1, a_curr_vec_in_AY_dqdPE1, a_curr_vec_in_AZ_dqdPE1, a_curr_vec_in_LX_dqdPE1, a_curr_vec_in_LY_dqdPE1, a_curr_vec_in_LZ_dqdPE1, a_curr_vec_in_AX_dqdPE2, a_curr_vec_in_AY_dqdPE2, a_curr_vec_in_AZ_dqdPE2, a_curr_vec_in_LX_dqdPE2, a_curr_vec_in_LY_dqdPE2, a_curr_vec_in_LZ_dqdPE2, a_curr_vec_in_AX_dqdPE3, a_curr_vec_in_AY_dqdPE3, a_curr_vec_in_AZ_dqdPE3, a_curr_vec_in_LX_dqdPE3, a_curr_vec_in_LY_dqdPE3, a_curr_vec_in_LZ_dqdPE3, a_curr_vec_in_AX_dqdPE4, a_curr_vec_in_AY_dqdPE4, a_curr_vec_in_AZ_dqdPE4, a_curr_vec_in_LX_dqdPE4, a_curr_vec_in_LY_dqdPE4, a_curr_vec_in_LZ_dqdPE4, a_curr_vec_in_AX_dqdPE5, a_curr_vec_in_AY_dqdPE5, a_curr_vec_in_AZ_dqdPE5, a_curr_vec_in_LX_dqdPE5, a_curr_vec_in_LY_dqdPE5, a_curr_vec_in_LZ_dqdPE5, a_curr_vec_in_AX_dqdPE6, a_curr_vec_in_AY_dqdPE6, a_curr_vec_in_AZ_dqdPE6, a_curr_vec_in_LX_dqdPE6, a_curr_vec_in_LY_dqdPE6, a_curr_vec_in_LZ_dqdPE6, a_curr_vec_in_AX_dqdPE7, a_curr_vec_in_AY_dqdPE7, a_curr_vec_in_AZ_dqdPE7, a_curr_vec_in_LX_dqdPE7, a_curr_vec_in_LY_dqdPE7, a_curr_vec_in_LZ_dqdPE7, v_prev_vec_in_AX_dqPE1, v_prev_vec_in_AY_dqPE1, v_prev_vec_in_AZ_dqPE1, v_prev_vec_in_LX_dqPE1, v_prev_vec_in_LY_dqPE1, v_prev_vec_in_LZ_dqPE1, v_prev_vec_in_AX_dqPE2, v_prev_vec_in_AY_dqPE2, v_prev_vec_in_AZ_dqPE2, v_prev_vec_in_LX_dqPE2, v_prev_vec_in_LY_dqPE2, v_prev_vec_in_LZ_dqPE2, v_prev_vec_in_AX_dqPE3, v_prev_vec_in_AY_dqPE3, v_prev_vec_in_AZ_dqPE3, v_prev_vec_in_LX_dqPE3, v_prev_vec_in_LY_dqPE3, v_prev_vec_in_LZ_dqPE3, v_prev_vec_in_AX_dqPE4, v_prev_vec_in_AY_dqPE4, v_prev_vec_in_AZ_dqPE4, v_prev_vec_in_LX_dqPE4, v_prev_vec_in_LY_dqPE4, v_prev_vec_in_LZ_dqPE4, v_prev_vec_in_AX_dqPE5, v_prev_vec_in_AY_dqPE5, v_prev_vec_in_AZ_dqPE5, v_prev_vec_in_LX_dqPE5, v_prev_vec_in_LY_dqPE5, v_prev_vec_in_LZ_dqPE5, v_prev_vec_in_AX_dqPE6, v_prev_vec_in_AY_dqPE6, v_prev_vec_in_AZ_dqPE6, v_prev_vec_in_LX_dqPE6, v_prev_vec_in_LY_dqPE6, v_prev_vec_in_LZ_dqPE6, v_prev_vec_in_AX_dqPE7, v_prev_vec_in_AY_dqPE7, v_prev_vec_in_AZ_dqPE7, v_prev_vec_in_LX_dqPE7, v_prev_vec_in_LY_dqPE7, v_prev_vec_in_LZ_dqPE7, a_prev_vec_in_AX_dqPE1, a_prev_vec_in_AY_dqPE1, a_prev_vec_in_AZ_dqPE1, a_prev_vec_in_LX_dqPE1, a_prev_vec_in_LY_dqPE1, a_prev_vec_in_LZ_dqPE1, a_prev_vec_in_AX_dqPE2, a_prev_vec_in_AY_dqPE2, a_prev_vec_in_AZ_dqPE2, a_prev_vec_in_LX_dqPE2, a_prev_vec_in_LY_dqPE2, a_prev_vec_in_LZ_dqPE2, a_prev_vec_in_AX_dqPE3, a_prev_vec_in_AY_dqPE3, a_prev_vec_in_AZ_dqPE3, a_prev_vec_in_LX_dqPE3, a_prev_vec_in_LY_dqPE3, a_prev_vec_in_LZ_dqPE3, a_prev_vec_in_AX_dqPE4, a_prev_vec_in_AY_dqPE4, a_prev_vec_in_AZ_dqPE4, a_prev_vec_in_LX_dqPE4, a_prev_vec_in_LY_dqPE4, a_prev_vec_in_LZ_dqPE4, a_prev_vec_in_AX_dqPE5, a_prev_vec_in_AY_dqPE5, a_prev_vec_in_AZ_dqPE5, a_prev_vec_in_LX_dqPE5, a_prev_vec_in_LY_dqPE5, a_prev_vec_in_LZ_dqPE5, a_prev_vec_in_AX_dqPE6, a_prev_vec_in_AY_dqPE6, a_prev_vec_in_AZ_dqPE6, a_prev_vec_in_LX_dqPE6, a_prev_vec_in_LY_dqPE6, a_prev_vec_in_LZ_dqPE6, a_prev_vec_in_AX_dqPE7, a_prev_vec_in_AY_dqPE7, a_prev_vec_in_AZ_dqPE7, a_prev_vec_in_LX_dqPE7, a_prev_vec_in_LY_dqPE7, a_prev_vec_in_LZ_dqPE7,
        dvdq_prev_vec_in_AX_dqPE1, dvdq_prev_vec_in_AY_dqPE1, dvdq_prev_vec_in_AZ_dqPE1, dvdq_prev_vec_in_LX_dqPE1, dvdq_prev_vec_in_LY_dqPE1, dvdq_prev_vec_in_LZ_dqPE1, dvdq_prev_vec_in_AX_dqPE2, dvdq_prev_vec_in_AY_dqPE2, dvdq_prev_vec_in_AZ_dqPE2, dvdq_prev_vec_in_LX_dqPE2, dvdq_prev_vec_in_LY_dqPE2, dvdq_prev_vec_in_LZ_dqPE2, dvdq_prev_vec_in_AX_dqPE3, dvdq_prev_vec_in_AY_dqPE3, dvdq_prev_vec_in_AZ_dqPE3, dvdq_prev_vec_in_LX_dqPE3, dvdq_prev_vec_in_LY_dqPE3, dvdq_prev_vec_in_LZ_dqPE3, dvdq_prev_vec_in_AX_dqPE4, dvdq_prev_vec_in_AY_dqPE4, dvdq_prev_vec_in_AZ_dqPE4, dvdq_prev_vec_in_LX_dqPE4, dvdq_prev_vec_in_LY_dqPE4, dvdq_prev_vec_in_LZ_dqPE4, dvdq_prev_vec_in_AX_dqPE5, dvdq_prev_vec_in_AY_dqPE5, dvdq_prev_vec_in_AZ_dqPE5, dvdq_prev_vec_in_LX_dqPE5, dvdq_prev_vec_in_LY_dqPE5, dvdq_prev_vec_in_LZ_dqPE5, dvdq_prev_vec_in_AX_dqPE6, dvdq_prev_vec_in_AY_dqPE6, dvdq_prev_vec_in_AZ_dqPE6, dvdq_prev_vec_in_LX_dqPE6, dvdq_prev_vec_in_LY_dqPE6, dvdq_prev_vec_in_LZ_dqPE6, dvdq_prev_vec_in_AX_dqPE7, dvdq_prev_vec_in_AY_dqPE7, dvdq_prev_vec_in_AZ_dqPE7, dvdq_prev_vec_in_LX_dqPE7, dvdq_prev_vec_in_LY_dqPE7, dvdq_prev_vec_in_LZ_dqPE7, dvdqd_prev_vec_in_AX_dqdPE1, dvdqd_prev_vec_in_AY_dqdPE1, dvdqd_prev_vec_in_AZ_dqdPE1, dvdqd_prev_vec_in_LX_dqdPE1, dvdqd_prev_vec_in_LY_dqdPE1, dvdqd_prev_vec_in_LZ_dqdPE1, dvdqd_prev_vec_in_AX_dqdPE2, dvdqd_prev_vec_in_AY_dqdPE2, dvdqd_prev_vec_in_AZ_dqdPE2, dvdqd_prev_vec_in_LX_dqdPE2, dvdqd_prev_vec_in_LY_dqdPE2, dvdqd_prev_vec_in_LZ_dqdPE2, dvdqd_prev_vec_in_AX_dqdPE3, dvdqd_prev_vec_in_AY_dqdPE3, dvdqd_prev_vec_in_AZ_dqdPE3, dvdqd_prev_vec_in_LX_dqdPE3, dvdqd_prev_vec_in_LY_dqdPE3, dvdqd_prev_vec_in_LZ_dqdPE3, dvdqd_prev_vec_in_AX_dqdPE4, dvdqd_prev_vec_in_AY_dqdPE4, dvdqd_prev_vec_in_AZ_dqdPE4, dvdqd_prev_vec_in_LX_dqdPE4, dvdqd_prev_vec_in_LY_dqdPE4, dvdqd_prev_vec_in_LZ_dqdPE4, dvdqd_prev_vec_in_AX_dqdPE5, dvdqd_prev_vec_in_AY_dqdPE5, dvdqd_prev_vec_in_AZ_dqdPE5, dvdqd_prev_vec_in_LX_dqdPE5, dvdqd_prev_vec_in_LY_dqdPE5, dvdqd_prev_vec_in_LZ_dqdPE5, dvdqd_prev_vec_in_AX_dqdPE6, dvdqd_prev_vec_in_AY_dqdPE6, dvdqd_prev_vec_in_AZ_dqdPE6, dvdqd_prev_vec_in_LX_dqdPE6, dvdqd_prev_vec_in_LY_dqdPE6, dvdqd_prev_vec_in_LZ_dqdPE6, dvdqd_prev_vec_in_AX_dqdPE7, dvdqd_prev_vec_in_AY_dqdPE7, dvdqd_prev_vec_in_AZ_dqdPE7, dvdqd_prev_vec_in_LX_dqdPE7, dvdqd_prev_vec_in_LY_dqdPE7, dvdqd_prev_vec_in_LZ_dqdPE7, dadq_prev_vec_in_AX_dqPE1, dadq_prev_vec_in_AY_dqPE1, dadq_prev_vec_in_AZ_dqPE1, dadq_prev_vec_in_LX_dqPE1, dadq_prev_vec_in_LY_dqPE1, dadq_prev_vec_in_LZ_dqPE1, dadq_prev_vec_in_AX_dqPE2, dadq_prev_vec_in_AY_dqPE2, dadq_prev_vec_in_AZ_dqPE2, dadq_prev_vec_in_LX_dqPE2, dadq_prev_vec_in_LY_dqPE2, dadq_prev_vec_in_LZ_dqPE2, dadq_prev_vec_in_AX_dqPE3, dadq_prev_vec_in_AY_dqPE3, dadq_prev_vec_in_AZ_dqPE3, dadq_prev_vec_in_LX_dqPE3, dadq_prev_vec_in_LY_dqPE3, dadq_prev_vec_in_LZ_dqPE3, dadq_prev_vec_in_AX_dqPE4, dadq_prev_vec_in_AY_dqPE4, dadq_prev_vec_in_AZ_dqPE4, dadq_prev_vec_in_LX_dqPE4, dadq_prev_vec_in_LY_dqPE4, dadq_prev_vec_in_LZ_dqPE4, dadq_prev_vec_in_AX_dqPE5, dadq_prev_vec_in_AY_dqPE5, dadq_prev_vec_in_AZ_dqPE5, dadq_prev_vec_in_LX_dqPE5, dadq_prev_vec_in_LY_dqPE5, dadq_prev_vec_in_LZ_dqPE5, dadq_prev_vec_in_AX_dqPE6, dadq_prev_vec_in_AY_dqPE6, dadq_prev_vec_in_AZ_dqPE6, dadq_prev_vec_in_LX_dqPE6, dadq_prev_vec_in_LY_dqPE6, dadq_prev_vec_in_LZ_dqPE6, dadq_prev_vec_in_AX_dqPE7, dadq_prev_vec_in_AY_dqPE7, dadq_prev_vec_in_AZ_dqPE7, dadq_prev_vec_in_LX_dqPE7, dadq_prev_vec_in_LY_dqPE7, dadq_prev_vec_in_LZ_dqPE7, dadqd_prev_vec_in_AX_dqdPE1, dadqd_prev_vec_in_AY_dqdPE1, dadqd_prev_vec_in_AZ_dqdPE1, dadqd_prev_vec_in_LX_dqdPE1, dadqd_prev_vec_in_LY_dqdPE1, dadqd_prev_vec_in_LZ_dqdPE1, dadqd_prev_vec_in_AX_dqdPE2, dadqd_prev_vec_in_AY_dqdPE2, dadqd_prev_vec_in_AZ_dqdPE2, dadqd_prev_vec_in_LX_dqdPE2, dadqd_prev_vec_in_LY_dqdPE2, dadqd_prev_vec_in_LZ_dqdPE2, dadqd_prev_vec_in_AX_dqdPE3, dadqd_prev_vec_in_AY_dqdPE3, dadqd_prev_vec_in_AZ_dqdPE3, dadqd_prev_vec_in_LX_dqdPE3, dadqd_prev_vec_in_LY_dqdPE3, dadqd_prev_vec_in_LZ_dqdPE3, dadqd_prev_vec_in_AX_dqdPE4, dadqd_prev_vec_in_AY_dqdPE4, dadqd_prev_vec_in_AZ_dqdPE4, dadqd_prev_vec_in_LX_dqdPE4, dadqd_prev_vec_in_LY_dqdPE4, dadqd_prev_vec_in_LZ_dqdPE4, dadqd_prev_vec_in_AX_dqdPE5, dadqd_prev_vec_in_AY_dqdPE5, dadqd_prev_vec_in_AZ_dqdPE5, dadqd_prev_vec_in_LX_dqdPE5, dadqd_prev_vec_in_LY_dqdPE5, dadqd_prev_vec_in_LZ_dqdPE5, dadqd_prev_vec_in_AX_dqdPE6, dadqd_prev_vec_in_AY_dqdPE6, dadqd_prev_vec_in_AZ_dqdPE6, dadqd_prev_vec_in_LX_dqdPE6, dadqd_prev_vec_in_LY_dqdPE6, dadqd_prev_vec_in_LZ_dqdPE6, dadqd_prev_vec_in_AX_dqdPE7, dadqd_prev_vec_in_AY_dqdPE7, dadqd_prev_vec_in_AZ_dqdPE7, dadqd_prev_vec_in_LX_dqdPE7, dadqd_prev_vec_in_LY_dqdPE7, dadqd_prev_vec_in_LZ_dqdPE7,
         output_ready,
        v_curr_vec_out_AX_rnea, v_curr_vec_out_AY_rnea, v_curr_vec_out_AZ_rnea, v_curr_vec_out_LX_rnea, v_curr_vec_out_LY_rnea, v_curr_vec_out_LZ_rnea, a_curr_vec_out_AX_rnea, a_curr_vec_out_AY_rnea, a_curr_vec_out_AZ_rnea, a_curr_vec_out_LX_rnea, a_curr_vec_out_LY_rnea, a_curr_vec_out_LZ_rnea, f_curr_vec_out_AX_rnea, f_curr_vec_out_AY_rnea, f_curr_vec_out_AZ_rnea, f_curr_vec_out_LX_rnea, f_curr_vec_out_LY_rnea, f_curr_vec_out_LZ_rnea,
        dfdq_curr_vec_out_AX_dqPE1, dfdq_curr_vec_out_AY_dqPE1, dfdq_curr_vec_out_AZ_dqPE1, dfdq_curr_vec_out_LX_dqPE1, dfdq_curr_vec_out_LY_dqPE1, dfdq_curr_vec_out_LZ_dqPE1, dfdq_curr_vec_out_AX_dqPE2, dfdq_curr_vec_out_AY_dqPE2, dfdq_curr_vec_out_AZ_dqPE2, dfdq_curr_vec_out_LX_dqPE2, dfdq_curr_vec_out_LY_dqPE2, dfdq_curr_vec_out_LZ_dqPE2, dfdq_curr_vec_out_AX_dqPE3, dfdq_curr_vec_out_AY_dqPE3, dfdq_curr_vec_out_AZ_dqPE3, dfdq_curr_vec_out_LX_dqPE3, dfdq_curr_vec_out_LY_dqPE3, dfdq_curr_vec_out_LZ_dqPE3, dfdq_curr_vec_out_AX_dqPE4, dfdq_curr_vec_out_AY_dqPE4, dfdq_curr_vec_out_AZ_dqPE4, dfdq_curr_vec_out_LX_dqPE4, dfdq_curr_vec_out_LY_dqPE4, dfdq_curr_vec_out_LZ_dqPE4, dfdq_curr_vec_out_AX_dqPE5, dfdq_curr_vec_out_AY_dqPE5, dfdq_curr_vec_out_AZ_dqPE5, dfdq_curr_vec_out_LX_dqPE5, dfdq_curr_vec_out_LY_dqPE5, dfdq_curr_vec_out_LZ_dqPE5, dfdq_curr_vec_out_AX_dqPE6, dfdq_curr_vec_out_AY_dqPE6, dfdq_curr_vec_out_AZ_dqPE6, dfdq_curr_vec_out_LX_dqPE6, dfdq_curr_vec_out_LY_dqPE6, dfdq_curr_vec_out_LZ_dqPE6, dfdq_curr_vec_out_AX_dqPE7, dfdq_curr_vec_out_AY_dqPE7, dfdq_curr_vec_out_AZ_dqPE7, dfdq_curr_vec_out_LX_dqPE7, dfdq_curr_vec_out_LY_dqPE7, dfdq_curr_vec_out_LZ_dqPE7, dfdqd_curr_vec_out_AX_dqdPE1, dfdqd_curr_vec_out_AY_dqdPE1, dfdqd_curr_vec_out_AZ_dqdPE1, dfdqd_curr_vec_out_LX_dqdPE1, dfdqd_curr_vec_out_LY_dqdPE1, dfdqd_curr_vec_out_LZ_dqdPE1, dfdqd_curr_vec_out_AX_dqdPE2, dfdqd_curr_vec_out_AY_dqdPE2, dfdqd_curr_vec_out_AZ_dqdPE2, dfdqd_curr_vec_out_LX_dqdPE2, dfdqd_curr_vec_out_LY_dqdPE2, dfdqd_curr_vec_out_LZ_dqdPE2, dfdqd_curr_vec_out_AX_dqdPE3, dfdqd_curr_vec_out_AY_dqdPE3, dfdqd_curr_vec_out_AZ_dqdPE3, dfdqd_curr_vec_out_LX_dqdPE3, dfdqd_curr_vec_out_LY_dqdPE3, dfdqd_curr_vec_out_LZ_dqdPE3, dfdqd_curr_vec_out_AX_dqdPE4, dfdqd_curr_vec_out_AY_dqdPE4, dfdqd_curr_vec_out_AZ_dqdPE4, dfdqd_curr_vec_out_LX_dqdPE4, dfdqd_curr_vec_out_LY_dqdPE4, dfdqd_curr_vec_out_LZ_dqdPE4, dfdqd_curr_vec_out_AX_dqdPE5, dfdqd_curr_vec_out_AY_dqdPE5, dfdqd_curr_vec_out_AZ_dqdPE5, dfdqd_curr_vec_out_LX_dqdPE5, dfdqd_curr_vec_out_LY_dqdPE5, dfdqd_curr_vec_out_LZ_dqdPE5, dfdqd_curr_vec_out_AX_dqdPE6, dfdqd_curr_vec_out_AY_dqdPE6, dfdqd_curr_vec_out_AZ_dqdPE6, dfdqd_curr_vec_out_LX_dqdPE6, dfdqd_curr_vec_out_LY_dqdPE6, dfdqd_curr_vec_out_LZ_dqdPE6, dfdqd_curr_vec_out_AX_dqdPE7, dfdqd_curr_vec_out_AY_dqdPE7, dfdqd_curr_vec_out_AZ_dqdPE7, dfdqd_curr_vec_out_LX_dqdPE7, dfdqd_curr_vec_out_LY_dqdPE7, dfdqd_curr_vec_out_LZ_dqdPE7,
        dvdq_curr_vec_out_AX_dqPE1, dvdq_curr_vec_out_AY_dqPE1, dvdq_curr_vec_out_AZ_dqPE1, dvdq_curr_vec_out_LX_dqPE1, dvdq_curr_vec_out_LY_dqPE1, dvdq_curr_vec_out_LZ_dqPE1, dvdq_curr_vec_out_AX_dqPE2, dvdq_curr_vec_out_AY_dqPE2, dvdq_curr_vec_out_AZ_dqPE2, dvdq_curr_vec_out_LX_dqPE2, dvdq_curr_vec_out_LY_dqPE2, dvdq_curr_vec_out_LZ_dqPE2, dvdq_curr_vec_out_AX_dqPE3, dvdq_curr_vec_out_AY_dqPE3, dvdq_curr_vec_out_AZ_dqPE3, dvdq_curr_vec_out_LX_dqPE3, dvdq_curr_vec_out_LY_dqPE3, dvdq_curr_vec_out_LZ_dqPE3, dvdq_curr_vec_out_AX_dqPE4, dvdq_curr_vec_out_AY_dqPE4, dvdq_curr_vec_out_AZ_dqPE4, dvdq_curr_vec_out_LX_dqPE4, dvdq_curr_vec_out_LY_dqPE4, dvdq_curr_vec_out_LZ_dqPE4, dvdq_curr_vec_out_AX_dqPE5, dvdq_curr_vec_out_AY_dqPE5, dvdq_curr_vec_out_AZ_dqPE5, dvdq_curr_vec_out_LX_dqPE5, dvdq_curr_vec_out_LY_dqPE5, dvdq_curr_vec_out_LZ_dqPE5, dvdq_curr_vec_out_AX_dqPE6, dvdq_curr_vec_out_AY_dqPE6, dvdq_curr_vec_out_AZ_dqPE6, dvdq_curr_vec_out_LX_dqPE6, dvdq_curr_vec_out_LY_dqPE6, dvdq_curr_vec_out_LZ_dqPE6, dvdq_curr_vec_out_AX_dqPE7, dvdq_curr_vec_out_AY_dqPE7, dvdq_curr_vec_out_AZ_dqPE7, dvdq_curr_vec_out_LX_dqPE7, dvdq_curr_vec_out_LY_dqPE7, dvdq_curr_vec_out_LZ_dqPE7, dvdqd_curr_vec_out_AX_dqdPE1, dvdqd_curr_vec_out_AY_dqdPE1, dvdqd_curr_vec_out_AZ_dqdPE1, dvdqd_curr_vec_out_LX_dqdPE1, dvdqd_curr_vec_out_LY_dqdPE1, dvdqd_curr_vec_out_LZ_dqdPE1, dvdqd_curr_vec_out_AX_dqdPE2, dvdqd_curr_vec_out_AY_dqdPE2, dvdqd_curr_vec_out_AZ_dqdPE2, dvdqd_curr_vec_out_LX_dqdPE2, dvdqd_curr_vec_out_LY_dqdPE2, dvdqd_curr_vec_out_LZ_dqdPE2, dvdqd_curr_vec_out_AX_dqdPE3, dvdqd_curr_vec_out_AY_dqdPE3, dvdqd_curr_vec_out_AZ_dqdPE3, dvdqd_curr_vec_out_LX_dqdPE3, dvdqd_curr_vec_out_LY_dqdPE3, dvdqd_curr_vec_out_LZ_dqdPE3, dvdqd_curr_vec_out_AX_dqdPE4, dvdqd_curr_vec_out_AY_dqdPE4, dvdqd_curr_vec_out_AZ_dqdPE4, dvdqd_curr_vec_out_LX_dqdPE4, dvdqd_curr_vec_out_LY_dqdPE4, dvdqd_curr_vec_out_LZ_dqdPE4, dvdqd_curr_vec_out_AX_dqdPE5, dvdqd_curr_vec_out_AY_dqdPE5, dvdqd_curr_vec_out_AZ_dqdPE5, dvdqd_curr_vec_out_LX_dqdPE5, dvdqd_curr_vec_out_LY_dqdPE5, dvdqd_curr_vec_out_LZ_dqdPE5, dvdqd_curr_vec_out_AX_dqdPE6, dvdqd_curr_vec_out_AY_dqdPE6, dvdqd_curr_vec_out_AZ_dqdPE6, dvdqd_curr_vec_out_LX_dqdPE6, dvdqd_curr_vec_out_LY_dqdPE6, dvdqd_curr_vec_out_LZ_dqdPE6, dvdqd_curr_vec_out_AX_dqdPE7, dvdqd_curr_vec_out_AY_dqdPE7, dvdqd_curr_vec_out_AZ_dqdPE7, dvdqd_curr_vec_out_LX_dqdPE7, dvdqd_curr_vec_out_LY_dqdPE7, dvdqd_curr_vec_out_LZ_dqdPE7, dadq_curr_vec_out_AX_dqPE1, dadq_curr_vec_out_AY_dqPE1, dadq_curr_vec_out_AZ_dqPE1, dadq_curr_vec_out_LX_dqPE1, dadq_curr_vec_out_LY_dqPE1, dadq_curr_vec_out_LZ_dqPE1, dadq_curr_vec_out_AX_dqPE2, dadq_curr_vec_out_AY_dqPE2, dadq_curr_vec_out_AZ_dqPE2, dadq_curr_vec_out_LX_dqPE2, dadq_curr_vec_out_LY_dqPE2, dadq_curr_vec_out_LZ_dqPE2, dadq_curr_vec_out_AX_dqPE3, dadq_curr_vec_out_AY_dqPE3, dadq_curr_vec_out_AZ_dqPE3, dadq_curr_vec_out_LX_dqPE3, dadq_curr_vec_out_LY_dqPE3, dadq_curr_vec_out_LZ_dqPE3, dadq_curr_vec_out_AX_dqPE4, dadq_curr_vec_out_AY_dqPE4, dadq_curr_vec_out_AZ_dqPE4, dadq_curr_vec_out_LX_dqPE4, dadq_curr_vec_out_LY_dqPE4, dadq_curr_vec_out_LZ_dqPE4, dadq_curr_vec_out_AX_dqPE5, dadq_curr_vec_out_AY_dqPE5, dadq_curr_vec_out_AZ_dqPE5, dadq_curr_vec_out_LX_dqPE5, dadq_curr_vec_out_LY_dqPE5, dadq_curr_vec_out_LZ_dqPE5, dadq_curr_vec_out_AX_dqPE6, dadq_curr_vec_out_AY_dqPE6, dadq_curr_vec_out_AZ_dqPE6, dadq_curr_vec_out_LX_dqPE6, dadq_curr_vec_out_LY_dqPE6, dadq_curr_vec_out_LZ_dqPE6, dadq_curr_vec_out_AX_dqPE7, dadq_curr_vec_out_AY_dqPE7, dadq_curr_vec_out_AZ_dqPE7, dadq_curr_vec_out_LX_dqPE7, dadq_curr_vec_out_LY_dqPE7, dadq_curr_vec_out_LZ_dqPE7, dadqd_curr_vec_out_AX_dqdPE1, dadqd_curr_vec_out_AY_dqdPE1, dadqd_curr_vec_out_AZ_dqdPE1, dadqd_curr_vec_out_LX_dqdPE1, dadqd_curr_vec_out_LY_dqdPE1, dadqd_curr_vec_out_LZ_dqdPE1, dadqd_curr_vec_out_AX_dqdPE2, dadqd_curr_vec_out_AY_dqdPE2, dadqd_curr_vec_out_AZ_dqdPE2, dadqd_curr_vec_out_LX_dqdPE2, dadqd_curr_vec_out_LY_dqdPE2, dadqd_curr_vec_out_LZ_dqdPE2, dadqd_curr_vec_out_AX_dqdPE3, dadqd_curr_vec_out_AY_dqdPE3, dadqd_curr_vec_out_AZ_dqdPE3, dadqd_curr_vec_out_LX_dqdPE3, dadqd_curr_vec_out_LY_dqdPE3, dadqd_curr_vec_out_LZ_dqdPE3, dadqd_curr_vec_out_AX_dqdPE4, dadqd_curr_vec_out_AY_dqdPE4, dadqd_curr_vec_out_AZ_dqdPE4, dadqd_curr_vec_out_LX_dqdPE4, dadqd_curr_vec_out_LY_dqdPE4, dadqd_curr_vec_out_LZ_dqdPE4, dadqd_curr_vec_out_AX_dqdPE5, dadqd_curr_vec_out_AY_dqdPE5, dadqd_curr_vec_out_AZ_dqdPE5, dadqd_curr_vec_out_LX_dqdPE5, dadqd_curr_vec_out_LY_dqdPE5, dadqd_curr_vec_out_LZ_dqdPE5, dadqd_curr_vec_out_AX_dqdPE6, dadqd_curr_vec_out_AY_dqdPE6, dadqd_curr_vec_out_AZ_dqdPE6, dadqd_curr_vec_out_LX_dqdPE6, dadqd_curr_vec_out_LY_dqdPE6, dadqd_curr_vec_out_LZ_dqdPE6, dadqd_curr_vec_out_AX_dqdPE7, dadqd_curr_vec_out_AY_dqdPE7, dadqd_curr_vec_out_AZ_dqdPE7, dadqd_curr_vec_out_LX_dqdPE7, dadqd_curr_vec_out_LY_dqdPE7, dadqd_curr_vec_out_LZ_dqdPE7
    );

endmodule
