Bit#(32) minv_block_in_R1_C1_dqdPE1 = 0;
Bit#(32) minv_block_in_R2_C1_dqdPE1 = 0;
Bit#(32) minv_block_in_R3_C1_dqdPE1 = 0;
Bit#(32) minv_block_in_R4_C1_dqdPE1 = 0;
Bit#(32) minv_block_in_R5_C1_dqdPE1 = 0;
Bit#(32) minv_block_in_R6_C1_dqdPE1 = 0;
Bit#(32) minv_block_in_R7_C1_dqdPE1 = 0;
Bit#(32) minv_block_in_R1_C2_dqdPE1 = 0;
Bit#(32) minv_block_in_R2_C2_dqdPE1 = 0;
Bit#(32) minv_block_in_R3_C2_dqdPE1 = 0;
Bit#(32) minv_block_in_R4_C2_dqdPE1 = 0;
Bit#(32) minv_block_in_R5_C2_dqdPE1 = 0;
Bit#(32) minv_block_in_R6_C2_dqdPE1 = 0;
Bit#(32) minv_block_in_R7_C2_dqdPE1 = 0;
Bit#(32) minv_block_in_R1_C3_dqdPE1 = 0;
Bit#(32) minv_block_in_R2_C3_dqdPE1 = 0;
Bit#(32) minv_block_in_R3_C3_dqdPE1 = 0;
Bit#(32) minv_block_in_R4_C3_dqdPE1 = 0;
Bit#(32) minv_block_in_R5_C3_dqdPE1 = 0;
Bit#(32) minv_block_in_R6_C3_dqdPE1 = 0;
Bit#(32) minv_block_in_R7_C3_dqdPE1 = 0;
Bit#(32) minv_block_in_R1_C4_dqdPE1 = 0;
Bit#(32) minv_block_in_R2_C4_dqdPE1 = 0;
Bit#(32) minv_block_in_R3_C4_dqdPE1 = 0;
Bit#(32) minv_block_in_R4_C4_dqdPE1 = 0;
Bit#(32) minv_block_in_R5_C4_dqdPE1 = 0;
Bit#(32) minv_block_in_R6_C4_dqdPE1 = 0;
Bit#(32) minv_block_in_R7_C4_dqdPE1 = 0;
Bit#(32) minv_block_in_R1_C5_dqdPE1 = 0;
Bit#(32) minv_block_in_R2_C5_dqdPE1 = 0;
Bit#(32) minv_block_in_R3_C5_dqdPE1 = 0;
Bit#(32) minv_block_in_R4_C5_dqdPE1 = 0;
Bit#(32) minv_block_in_R5_C5_dqdPE1 = 0;
Bit#(32) minv_block_in_R6_C5_dqdPE1 = 0;
Bit#(32) minv_block_in_R7_C5_dqdPE1 = 0;
Bit#(32) minv_block_in_R1_C6_dqdPE1 = 0;
Bit#(32) minv_block_in_R2_C6_dqdPE1 = 0;
Bit#(32) minv_block_in_R3_C6_dqdPE1 = 0;
Bit#(32) minv_block_in_R4_C6_dqdPE1 = 0;
Bit#(32) minv_block_in_R5_C6_dqdPE1 = 0;
Bit#(32) minv_block_in_R6_C6_dqdPE1 = 0;
Bit#(32) minv_block_in_R7_C6_dqdPE1 = 0;
Bit#(32) minv_block_in_R1_C7_dqdPE1 = 0;
Bit#(32) minv_block_in_R2_C7_dqdPE1 = 0;
Bit#(32) minv_block_in_R3_C7_dqdPE1 = 0;
Bit#(32) minv_block_in_R4_C7_dqdPE1 = 0;
Bit#(32) minv_block_in_R5_C7_dqdPE1 = 0;
Bit#(32) minv_block_in_R6_C7_dqdPE1 = 0;
Bit#(32) minv_block_in_R7_C7_dqdPE1 = 0;
Bit#(32) minv_block_in_R1_C1_dqdPE2 = 0;
Bit#(32) minv_block_in_R2_C1_dqdPE2 = 0;
Bit#(32) minv_block_in_R3_C1_dqdPE2 = 0;
Bit#(32) minv_block_in_R4_C1_dqdPE2 = 0;
Bit#(32) minv_block_in_R5_C1_dqdPE2 = 0;
Bit#(32) minv_block_in_R6_C1_dqdPE2 = 0;
Bit#(32) minv_block_in_R7_C1_dqdPE2 = 0;
Bit#(32) minv_block_in_R1_C2_dqdPE2 = 0;
Bit#(32) minv_block_in_R2_C2_dqdPE2 = 0;
Bit#(32) minv_block_in_R3_C2_dqdPE2 = 0;
Bit#(32) minv_block_in_R4_C2_dqdPE2 = 0;
Bit#(32) minv_block_in_R5_C2_dqdPE2 = 0;
Bit#(32) minv_block_in_R6_C2_dqdPE2 = 0;
Bit#(32) minv_block_in_R7_C2_dqdPE2 = 0;
Bit#(32) minv_block_in_R1_C3_dqdPE2 = 0;
Bit#(32) minv_block_in_R2_C3_dqdPE2 = 0;
Bit#(32) minv_block_in_R3_C3_dqdPE2 = 0;
Bit#(32) minv_block_in_R4_C3_dqdPE2 = 0;
Bit#(32) minv_block_in_R5_C3_dqdPE2 = 0;
Bit#(32) minv_block_in_R6_C3_dqdPE2 = 0;
Bit#(32) minv_block_in_R7_C3_dqdPE2 = 0;
Bit#(32) minv_block_in_R1_C4_dqdPE2 = 0;
Bit#(32) minv_block_in_R2_C4_dqdPE2 = 0;
Bit#(32) minv_block_in_R3_C4_dqdPE2 = 0;
Bit#(32) minv_block_in_R4_C4_dqdPE2 = 0;
Bit#(32) minv_block_in_R5_C4_dqdPE2 = 0;
Bit#(32) minv_block_in_R6_C4_dqdPE2 = 0;
Bit#(32) minv_block_in_R7_C4_dqdPE2 = 0;
Bit#(32) minv_block_in_R1_C5_dqdPE2 = 0;
Bit#(32) minv_block_in_R2_C5_dqdPE2 = 0;
Bit#(32) minv_block_in_R3_C5_dqdPE2 = 0;
Bit#(32) minv_block_in_R4_C5_dqdPE2 = 0;
Bit#(32) minv_block_in_R5_C5_dqdPE2 = 0;
Bit#(32) minv_block_in_R6_C5_dqdPE2 = 0;
Bit#(32) minv_block_in_R7_C5_dqdPE2 = 0;
Bit#(32) minv_block_in_R1_C6_dqdPE2 = 0;
Bit#(32) minv_block_in_R2_C6_dqdPE2 = 0;
Bit#(32) minv_block_in_R3_C6_dqdPE2 = 0;
Bit#(32) minv_block_in_R4_C6_dqdPE2 = 0;
Bit#(32) minv_block_in_R5_C6_dqdPE2 = 0;
Bit#(32) minv_block_in_R6_C6_dqdPE2 = 0;
Bit#(32) minv_block_in_R7_C6_dqdPE2 = 0;
Bit#(32) minv_block_in_R1_C7_dqdPE2 = 0;
Bit#(32) minv_block_in_R2_C7_dqdPE2 = 0;
Bit#(32) minv_block_in_R3_C7_dqdPE2 = 0;
Bit#(32) minv_block_in_R4_C7_dqdPE2 = 0;
Bit#(32) minv_block_in_R5_C7_dqdPE2 = 0;
Bit#(32) minv_block_in_R6_C7_dqdPE2 = 0;
Bit#(32) minv_block_in_R7_C7_dqdPE2 = 0;
Bit#(32) minv_block_in_R1_C1_dqdPE3 = 0;
Bit#(32) minv_block_in_R2_C1_dqdPE3 = 0;
Bit#(32) minv_block_in_R3_C1_dqdPE3 = 0;
Bit#(32) minv_block_in_R4_C1_dqdPE3 = 0;
Bit#(32) minv_block_in_R5_C1_dqdPE3 = 0;
Bit#(32) minv_block_in_R6_C1_dqdPE3 = 0;
Bit#(32) minv_block_in_R7_C1_dqdPE3 = 0;
Bit#(32) minv_block_in_R1_C2_dqdPE3 = 0;
Bit#(32) minv_block_in_R2_C2_dqdPE3 = 0;
Bit#(32) minv_block_in_R3_C2_dqdPE3 = 0;
Bit#(32) minv_block_in_R4_C2_dqdPE3 = 0;
Bit#(32) minv_block_in_R5_C2_dqdPE3 = 0;
Bit#(32) minv_block_in_R6_C2_dqdPE3 = 0;
Bit#(32) minv_block_in_R7_C2_dqdPE3 = 0;
Bit#(32) minv_block_in_R1_C3_dqdPE3 = 0;
Bit#(32) minv_block_in_R2_C3_dqdPE3 = 0;
Bit#(32) minv_block_in_R3_C3_dqdPE3 = 0;
Bit#(32) minv_block_in_R4_C3_dqdPE3 = 0;
Bit#(32) minv_block_in_R5_C3_dqdPE3 = 0;
Bit#(32) minv_block_in_R6_C3_dqdPE3 = 0;
Bit#(32) minv_block_in_R7_C3_dqdPE3 = 0;
Bit#(32) minv_block_in_R1_C4_dqdPE3 = 0;
Bit#(32) minv_block_in_R2_C4_dqdPE3 = 0;
Bit#(32) minv_block_in_R3_C4_dqdPE3 = 0;
Bit#(32) minv_block_in_R4_C4_dqdPE3 = 0;
Bit#(32) minv_block_in_R5_C4_dqdPE3 = 0;
Bit#(32) minv_block_in_R6_C4_dqdPE3 = 0;
Bit#(32) minv_block_in_R7_C4_dqdPE3 = 0;
Bit#(32) minv_block_in_R1_C5_dqdPE3 = 0;
Bit#(32) minv_block_in_R2_C5_dqdPE3 = 0;
Bit#(32) minv_block_in_R3_C5_dqdPE3 = 0;
Bit#(32) minv_block_in_R4_C5_dqdPE3 = 0;
Bit#(32) minv_block_in_R5_C5_dqdPE3 = 0;
Bit#(32) minv_block_in_R6_C5_dqdPE3 = 0;
Bit#(32) minv_block_in_R7_C5_dqdPE3 = 0;
Bit#(32) minv_block_in_R1_C6_dqdPE3 = 0;
Bit#(32) minv_block_in_R2_C6_dqdPE3 = 0;
Bit#(32) minv_block_in_R3_C6_dqdPE3 = 0;
Bit#(32) minv_block_in_R4_C6_dqdPE3 = 0;
Bit#(32) minv_block_in_R5_C6_dqdPE3 = 0;
Bit#(32) minv_block_in_R6_C6_dqdPE3 = 0;
Bit#(32) minv_block_in_R7_C6_dqdPE3 = 0;
Bit#(32) minv_block_in_R1_C7_dqdPE3 = 0;
Bit#(32) minv_block_in_R2_C7_dqdPE3 = 0;
Bit#(32) minv_block_in_R3_C7_dqdPE3 = 0;
Bit#(32) minv_block_in_R4_C7_dqdPE3 = 0;
Bit#(32) minv_block_in_R5_C7_dqdPE3 = 0;
Bit#(32) minv_block_in_R6_C7_dqdPE3 = 0;
Bit#(32) minv_block_in_R7_C7_dqdPE3 = 0;
Bit#(32) minv_block_in_R1_C1_dqdPE4 = 0;
Bit#(32) minv_block_in_R2_C1_dqdPE4 = 0;
Bit#(32) minv_block_in_R3_C1_dqdPE4 = 0;
Bit#(32) minv_block_in_R4_C1_dqdPE4 = 0;
Bit#(32) minv_block_in_R5_C1_dqdPE4 = 0;
Bit#(32) minv_block_in_R6_C1_dqdPE4 = 0;
Bit#(32) minv_block_in_R7_C1_dqdPE4 = 0;
Bit#(32) minv_block_in_R1_C2_dqdPE4 = 0;
Bit#(32) minv_block_in_R2_C2_dqdPE4 = 0;
Bit#(32) minv_block_in_R3_C2_dqdPE4 = 0;
Bit#(32) minv_block_in_R4_C2_dqdPE4 = 0;
Bit#(32) minv_block_in_R5_C2_dqdPE4 = 0;
Bit#(32) minv_block_in_R6_C2_dqdPE4 = 0;
Bit#(32) minv_block_in_R7_C2_dqdPE4 = 0;
Bit#(32) minv_block_in_R1_C3_dqdPE4 = 0;
Bit#(32) minv_block_in_R2_C3_dqdPE4 = 0;
Bit#(32) minv_block_in_R3_C3_dqdPE4 = 0;
Bit#(32) minv_block_in_R4_C3_dqdPE4 = 0;
Bit#(32) minv_block_in_R5_C3_dqdPE4 = 0;
Bit#(32) minv_block_in_R6_C3_dqdPE4 = 0;
Bit#(32) minv_block_in_R7_C3_dqdPE4 = 0;
Bit#(32) minv_block_in_R1_C4_dqdPE4 = 0;
Bit#(32) minv_block_in_R2_C4_dqdPE4 = 0;
Bit#(32) minv_block_in_R3_C4_dqdPE4 = 0;
Bit#(32) minv_block_in_R4_C4_dqdPE4 = 0;
Bit#(32) minv_block_in_R5_C4_dqdPE4 = 0;
Bit#(32) minv_block_in_R6_C4_dqdPE4 = 0;
Bit#(32) minv_block_in_R7_C4_dqdPE4 = 0;
Bit#(32) minv_block_in_R1_C5_dqdPE4 = 0;
Bit#(32) minv_block_in_R2_C5_dqdPE4 = 0;
Bit#(32) minv_block_in_R3_C5_dqdPE4 = 0;
Bit#(32) minv_block_in_R4_C5_dqdPE4 = 0;
Bit#(32) minv_block_in_R5_C5_dqdPE4 = 0;
Bit#(32) minv_block_in_R6_C5_dqdPE4 = 0;
Bit#(32) minv_block_in_R7_C5_dqdPE4 = 0;
Bit#(32) minv_block_in_R1_C6_dqdPE4 = 0;
Bit#(32) minv_block_in_R2_C6_dqdPE4 = 0;
Bit#(32) minv_block_in_R3_C6_dqdPE4 = 0;
Bit#(32) minv_block_in_R4_C6_dqdPE4 = 0;
Bit#(32) minv_block_in_R5_C6_dqdPE4 = 0;
Bit#(32) minv_block_in_R6_C6_dqdPE4 = 0;
Bit#(32) minv_block_in_R7_C6_dqdPE4 = 0;
Bit#(32) minv_block_in_R1_C7_dqdPE4 = 0;
Bit#(32) minv_block_in_R2_C7_dqdPE4 = 0;
Bit#(32) minv_block_in_R3_C7_dqdPE4 = 0;
Bit#(32) minv_block_in_R4_C7_dqdPE4 = 0;
Bit#(32) minv_block_in_R5_C7_dqdPE4 = 0;
Bit#(32) minv_block_in_R6_C7_dqdPE4 = 0;
Bit#(32) minv_block_in_R7_C7_dqdPE4 = 0;
Bit#(32) minv_block_in_R1_C1_dqdPE5 = 0;
Bit#(32) minv_block_in_R2_C1_dqdPE5 = 0;
Bit#(32) minv_block_in_R3_C1_dqdPE5 = 0;
Bit#(32) minv_block_in_R4_C1_dqdPE5 = 0;
Bit#(32) minv_block_in_R5_C1_dqdPE5 = 0;
Bit#(32) minv_block_in_R6_C1_dqdPE5 = 0;
Bit#(32) minv_block_in_R7_C1_dqdPE5 = 0;
Bit#(32) minv_block_in_R1_C2_dqdPE5 = 0;
Bit#(32) minv_block_in_R2_C2_dqdPE5 = 0;
Bit#(32) minv_block_in_R3_C2_dqdPE5 = 0;
Bit#(32) minv_block_in_R4_C2_dqdPE5 = 0;
Bit#(32) minv_block_in_R5_C2_dqdPE5 = 0;
Bit#(32) minv_block_in_R6_C2_dqdPE5 = 0;
Bit#(32) minv_block_in_R7_C2_dqdPE5 = 0;
Bit#(32) minv_block_in_R1_C3_dqdPE5 = 0;
Bit#(32) minv_block_in_R2_C3_dqdPE5 = 0;
Bit#(32) minv_block_in_R3_C3_dqdPE5 = 0;
Bit#(32) minv_block_in_R4_C3_dqdPE5 = 0;
Bit#(32) minv_block_in_R5_C3_dqdPE5 = 0;
Bit#(32) minv_block_in_R6_C3_dqdPE5 = 0;
Bit#(32) minv_block_in_R7_C3_dqdPE5 = 0;
Bit#(32) minv_block_in_R1_C4_dqdPE5 = 0;
Bit#(32) minv_block_in_R2_C4_dqdPE5 = 0;
Bit#(32) minv_block_in_R3_C4_dqdPE5 = 0;
Bit#(32) minv_block_in_R4_C4_dqdPE5 = 0;
Bit#(32) minv_block_in_R5_C4_dqdPE5 = 0;
Bit#(32) minv_block_in_R6_C4_dqdPE5 = 0;
Bit#(32) minv_block_in_R7_C4_dqdPE5 = 0;
Bit#(32) minv_block_in_R1_C5_dqdPE5 = 0;
Bit#(32) minv_block_in_R2_C5_dqdPE5 = 0;
Bit#(32) minv_block_in_R3_C5_dqdPE5 = 0;
Bit#(32) minv_block_in_R4_C5_dqdPE5 = 0;
Bit#(32) minv_block_in_R5_C5_dqdPE5 = 0;
Bit#(32) minv_block_in_R6_C5_dqdPE5 = 0;
Bit#(32) minv_block_in_R7_C5_dqdPE5 = 0;
Bit#(32) minv_block_in_R1_C6_dqdPE5 = 0;
Bit#(32) minv_block_in_R2_C6_dqdPE5 = 0;
Bit#(32) minv_block_in_R3_C6_dqdPE5 = 0;
Bit#(32) minv_block_in_R4_C6_dqdPE5 = 0;
Bit#(32) minv_block_in_R5_C6_dqdPE5 = 0;
Bit#(32) minv_block_in_R6_C6_dqdPE5 = 0;
Bit#(32) minv_block_in_R7_C6_dqdPE5 = 0;
Bit#(32) minv_block_in_R1_C7_dqdPE5 = 0;
Bit#(32) minv_block_in_R2_C7_dqdPE5 = 0;
Bit#(32) minv_block_in_R3_C7_dqdPE5 = 0;
Bit#(32) minv_block_in_R4_C7_dqdPE5 = 0;
Bit#(32) minv_block_in_R5_C7_dqdPE5 = 0;
Bit#(32) minv_block_in_R6_C7_dqdPE5 = 0;
Bit#(32) minv_block_in_R7_C7_dqdPE5 = 0;
Bit#(32) minv_block_in_R1_C1_dqdPE6 = 0;
Bit#(32) minv_block_in_R2_C1_dqdPE6 = 0;
Bit#(32) minv_block_in_R3_C1_dqdPE6 = 0;
Bit#(32) minv_block_in_R4_C1_dqdPE6 = 0;
Bit#(32) minv_block_in_R5_C1_dqdPE6 = 0;
Bit#(32) minv_block_in_R6_C1_dqdPE6 = 0;
Bit#(32) minv_block_in_R7_C1_dqdPE6 = 0;
Bit#(32) minv_block_in_R1_C2_dqdPE6 = 0;
Bit#(32) minv_block_in_R2_C2_dqdPE6 = 0;
Bit#(32) minv_block_in_R3_C2_dqdPE6 = 0;
Bit#(32) minv_block_in_R4_C2_dqdPE6 = 0;
Bit#(32) minv_block_in_R5_C2_dqdPE6 = 0;
Bit#(32) minv_block_in_R6_C2_dqdPE6 = 0;
Bit#(32) minv_block_in_R7_C2_dqdPE6 = 0;
Bit#(32) minv_block_in_R1_C3_dqdPE6 = 0;
Bit#(32) minv_block_in_R2_C3_dqdPE6 = 0;
Bit#(32) minv_block_in_R3_C3_dqdPE6 = 0;
Bit#(32) minv_block_in_R4_C3_dqdPE6 = 0;
Bit#(32) minv_block_in_R5_C3_dqdPE6 = 0;
Bit#(32) minv_block_in_R6_C3_dqdPE6 = 0;
Bit#(32) minv_block_in_R7_C3_dqdPE6 = 0;
Bit#(32) minv_block_in_R1_C4_dqdPE6 = 0;
Bit#(32) minv_block_in_R2_C4_dqdPE6 = 0;
Bit#(32) minv_block_in_R3_C4_dqdPE6 = 0;
Bit#(32) minv_block_in_R4_C4_dqdPE6 = 0;
Bit#(32) minv_block_in_R5_C4_dqdPE6 = 0;
Bit#(32) minv_block_in_R6_C4_dqdPE6 = 0;
Bit#(32) minv_block_in_R7_C4_dqdPE6 = 0;
Bit#(32) minv_block_in_R1_C5_dqdPE6 = 0;
Bit#(32) minv_block_in_R2_C5_dqdPE6 = 0;
Bit#(32) minv_block_in_R3_C5_dqdPE6 = 0;
Bit#(32) minv_block_in_R4_C5_dqdPE6 = 0;
Bit#(32) minv_block_in_R5_C5_dqdPE6 = 0;
Bit#(32) minv_block_in_R6_C5_dqdPE6 = 0;
Bit#(32) minv_block_in_R7_C5_dqdPE6 = 0;
Bit#(32) minv_block_in_R1_C6_dqdPE6 = 0;
Bit#(32) minv_block_in_R2_C6_dqdPE6 = 0;
Bit#(32) minv_block_in_R3_C6_dqdPE6 = 0;
Bit#(32) minv_block_in_R4_C6_dqdPE6 = 0;
Bit#(32) minv_block_in_R5_C6_dqdPE6 = 0;
Bit#(32) minv_block_in_R6_C6_dqdPE6 = 0;
Bit#(32) minv_block_in_R7_C6_dqdPE6 = 0;
Bit#(32) minv_block_in_R1_C7_dqdPE6 = 0;
Bit#(32) minv_block_in_R2_C7_dqdPE6 = 0;
Bit#(32) minv_block_in_R3_C7_dqdPE6 = 0;
Bit#(32) minv_block_in_R4_C7_dqdPE6 = 0;
Bit#(32) minv_block_in_R5_C7_dqdPE6 = 0;
Bit#(32) minv_block_in_R6_C7_dqdPE6 = 0;
Bit#(32) minv_block_in_R7_C7_dqdPE6 = 0;
Bit#(32) minv_block_in_R1_C1_dqdPE7 = 0;
Bit#(32) minv_block_in_R2_C1_dqdPE7 = 0;
Bit#(32) minv_block_in_R3_C1_dqdPE7 = 0;
Bit#(32) minv_block_in_R4_C1_dqdPE7 = 0;
Bit#(32) minv_block_in_R5_C1_dqdPE7 = 0;
Bit#(32) minv_block_in_R6_C1_dqdPE7 = 0;
Bit#(32) minv_block_in_R7_C1_dqdPE7 = 0;
Bit#(32) minv_block_in_R1_C2_dqdPE7 = 0;
Bit#(32) minv_block_in_R2_C2_dqdPE7 = 0;
Bit#(32) minv_block_in_R3_C2_dqdPE7 = 0;
Bit#(32) minv_block_in_R4_C2_dqdPE7 = 0;
Bit#(32) minv_block_in_R5_C2_dqdPE7 = 0;
Bit#(32) minv_block_in_R6_C2_dqdPE7 = 0;
Bit#(32) minv_block_in_R7_C2_dqdPE7 = 0;
Bit#(32) minv_block_in_R1_C3_dqdPE7 = 0;
Bit#(32) minv_block_in_R2_C3_dqdPE7 = 0;
Bit#(32) minv_block_in_R3_C3_dqdPE7 = 0;
Bit#(32) minv_block_in_R4_C3_dqdPE7 = 0;
Bit#(32) minv_block_in_R5_C3_dqdPE7 = 0;
Bit#(32) minv_block_in_R6_C3_dqdPE7 = 0;
Bit#(32) minv_block_in_R7_C3_dqdPE7 = 0;
Bit#(32) minv_block_in_R1_C4_dqdPE7 = 0;
Bit#(32) minv_block_in_R2_C4_dqdPE7 = 0;
Bit#(32) minv_block_in_R3_C4_dqdPE7 = 0;
Bit#(32) minv_block_in_R4_C4_dqdPE7 = 0;
Bit#(32) minv_block_in_R5_C4_dqdPE7 = 0;
Bit#(32) minv_block_in_R6_C4_dqdPE7 = 0;
Bit#(32) minv_block_in_R7_C4_dqdPE7 = 0;
Bit#(32) minv_block_in_R1_C5_dqdPE7 = 0;
Bit#(32) minv_block_in_R2_C5_dqdPE7 = 0;
Bit#(32) minv_block_in_R3_C5_dqdPE7 = 0;
Bit#(32) minv_block_in_R4_C5_dqdPE7 = 0;
Bit#(32) minv_block_in_R5_C5_dqdPE7 = 0;
Bit#(32) minv_block_in_R6_C5_dqdPE7 = 0;
Bit#(32) minv_block_in_R7_C5_dqdPE7 = 0;
Bit#(32) minv_block_in_R1_C6_dqdPE7 = 0;
Bit#(32) minv_block_in_R2_C6_dqdPE7 = 0;
Bit#(32) minv_block_in_R3_C6_dqdPE7 = 0;
Bit#(32) minv_block_in_R4_C6_dqdPE7 = 0;
Bit#(32) minv_block_in_R5_C6_dqdPE7 = 0;
Bit#(32) minv_block_in_R6_C6_dqdPE7 = 0;
Bit#(32) minv_block_in_R7_C6_dqdPE7 = 0;
Bit#(32) minv_block_in_R1_C7_dqdPE7 = 0;
Bit#(32) minv_block_in_R2_C7_dqdPE7 = 0;
Bit#(32) minv_block_in_R3_C7_dqdPE7 = 0;
Bit#(32) minv_block_in_R4_C7_dqdPE7 = 0;
Bit#(32) minv_block_in_R5_C7_dqdPE7 = 0;
Bit#(32) minv_block_in_R6_C7_dqdPE7 = 0;
Bit#(32) minv_block_in_R7_C7_dqdPE7 = 0;

Bit#(32) dtau_vec_in_R1_dqdPE1 = 0;
Bit#(32) dtau_vec_in_R2_dqdPE1 = 0;
Bit#(32) dtau_vec_in_R3_dqdPE1 = 0;
Bit#(32) dtau_vec_in_R4_dqdPE1 = 0;
Bit#(32) dtau_vec_in_R5_dqdPE1 = 0;
Bit#(32) dtau_vec_in_R6_dqdPE1 = 0;
Bit#(32) dtau_vec_in_R7_dqdPE1 = 0;
Bit#(32) dtau_vec_in_R1_dqdPE2 = 0;
Bit#(32) dtau_vec_in_R2_dqdPE2 = 0;
Bit#(32) dtau_vec_in_R3_dqdPE2 = 0;
Bit#(32) dtau_vec_in_R4_dqdPE2 = 0;
Bit#(32) dtau_vec_in_R5_dqdPE2 = 0;
Bit#(32) dtau_vec_in_R6_dqdPE2 = 0;
Bit#(32) dtau_vec_in_R7_dqdPE2 = 0;
Bit#(32) dtau_vec_in_R1_dqdPE3 = 0;
Bit#(32) dtau_vec_in_R2_dqdPE3 = 0;
Bit#(32) dtau_vec_in_R3_dqdPE3 = 0;
Bit#(32) dtau_vec_in_R4_dqdPE3 = 0;
Bit#(32) dtau_vec_in_R5_dqdPE3 = 0;
Bit#(32) dtau_vec_in_R6_dqdPE3 = 0;
Bit#(32) dtau_vec_in_R7_dqdPE3 = 0;
Bit#(32) dtau_vec_in_R1_dqdPE4 = 0;
Bit#(32) dtau_vec_in_R2_dqdPE4 = 0;
Bit#(32) dtau_vec_in_R3_dqdPE4 = 0;
Bit#(32) dtau_vec_in_R4_dqdPE4 = 0;
Bit#(32) dtau_vec_in_R5_dqdPE4 = 0;
Bit#(32) dtau_vec_in_R6_dqdPE4 = 0;
Bit#(32) dtau_vec_in_R7_dqdPE4 = 0;
Bit#(32) dtau_vec_in_R1_dqdPE5 = 0;
Bit#(32) dtau_vec_in_R2_dqdPE5 = 0;
Bit#(32) dtau_vec_in_R3_dqdPE5 = 0;
Bit#(32) dtau_vec_in_R4_dqdPE5 = 0;
Bit#(32) dtau_vec_in_R5_dqdPE5 = 0;
Bit#(32) dtau_vec_in_R6_dqdPE5 = 0;
Bit#(32) dtau_vec_in_R7_dqdPE5 = 0;
Bit#(32) dtau_vec_in_R1_dqdPE6 = 0;
Bit#(32) dtau_vec_in_R2_dqdPE6 = 0;
Bit#(32) dtau_vec_in_R3_dqdPE6 = 0;
Bit#(32) dtau_vec_in_R4_dqdPE6 = 0;
Bit#(32) dtau_vec_in_R5_dqdPE6 = 0;
Bit#(32) dtau_vec_in_R6_dqdPE6 = 0;
Bit#(32) dtau_vec_in_R7_dqdPE6 = 0;
Bit#(32) dtau_vec_in_R1_dqdPE7 = 0;
Bit#(32) dtau_vec_in_R2_dqdPE7 = 0;
Bit#(32) dtau_vec_in_R3_dqdPE7 = 0;
Bit#(32) dtau_vec_in_R4_dqdPE7 = 0;
Bit#(32) dtau_vec_in_R5_dqdPE7 = 0;
Bit#(32) dtau_vec_in_R6_dqdPE7 = 0;
Bit#(32) dtau_vec_in_R7_dqdPE7 = 0;

case (idx_block_minv_feed_dtau)

    0: begin
        minv_block_in_R1_C1_dqdPE1 = minv[0][0];
        minv_block_in_R2_C1_dqdPE1 = minv[1][0];
        minv_block_in_R3_C1_dqdPE1 = minv[2][0];
        minv_block_in_R4_C1_dqdPE1 = minv[3][0];
        minv_block_in_R5_C1_dqdPE1 = minv[4][0];
        minv_block_in_R6_C1_dqdPE1 = minv[5][0];
        minv_block_in_R7_C1_dqdPE1 = minv[6][0];

        minv_block_in_R1_C2_dqdPE1 = minv[0][1];
        minv_block_in_R2_C2_dqdPE1 = minv[1][1];
        minv_block_in_R3_C2_dqdPE1 = minv[2][1];
        minv_block_in_R4_C2_dqdPE1 = minv[3][1];
        minv_block_in_R5_C2_dqdPE1 = minv[4][1];
        minv_block_in_R6_C2_dqdPE1 = minv[5][1];
        minv_block_in_R7_C2_dqdPE1 = minv[6][1];

        minv_block_in_R1_C3_dqdPE1 = minv[0][2];
        minv_block_in_R2_C3_dqdPE1 = minv[1][2];
        minv_block_in_R3_C3_dqdPE1 = minv[2][2];
        minv_block_in_R4_C3_dqdPE1 = minv[3][2];
        minv_block_in_R5_C3_dqdPE1 = minv[4][2];
        minv_block_in_R6_C3_dqdPE1 = minv[5][2];
        minv_block_in_R7_C3_dqdPE1 = minv[6][2];

        minv_block_in_R1_C4_dqdPE1 = minv[0][3];
        minv_block_in_R2_C4_dqdPE1 = minv[1][3];
        minv_block_in_R3_C4_dqdPE1 = minv[2][3];
        minv_block_in_R4_C4_dqdPE1 = minv[3][3];
        minv_block_in_R5_C4_dqdPE1 = minv[4][3];
        minv_block_in_R6_C4_dqdPE1 = minv[5][3];
        minv_block_in_R7_C4_dqdPE1 = minv[6][3];

        minv_block_in_R1_C5_dqdPE1 = minv[0][4];
        minv_block_in_R2_C5_dqdPE1 = minv[1][4];
        minv_block_in_R3_C5_dqdPE1 = minv[2][4];
        minv_block_in_R4_C5_dqdPE1 = minv[3][4];
        minv_block_in_R5_C5_dqdPE1 = minv[4][4];
        minv_block_in_R6_C5_dqdPE1 = minv[5][4];
        minv_block_in_R7_C5_dqdPE1 = minv[6][4];

        minv_block_in_R1_C6_dqdPE1 = minv[0][5];
        minv_block_in_R2_C6_dqdPE1 = minv[1][5];
        minv_block_in_R3_C6_dqdPE1 = minv[2][5];
        minv_block_in_R4_C6_dqdPE1 = minv[3][5];
        minv_block_in_R5_C6_dqdPE1 = minv[4][5];
        minv_block_in_R6_C6_dqdPE1 = minv[5][5];
        minv_block_in_R7_C6_dqdPE1 = minv[6][5];

        minv_block_in_R1_C7_dqdPE1 = minv[0][6];
        minv_block_in_R2_C7_dqdPE1 = minv[1][6];
        minv_block_in_R3_C7_dqdPE1 = minv[2][6];
        minv_block_in_R4_C7_dqdPE1 = minv[3][6];
        minv_block_in_R5_C7_dqdPE1 = minv[4][6];
        minv_block_in_R6_C7_dqdPE1 = minv[5][6];
        minv_block_in_R7_C7_dqdPE1 = minv[6][6];

        minv_block_in_R1_C1_dqdPE2 = minv[0][0];
        minv_block_in_R2_C1_dqdPE2 = minv[1][0];
        minv_block_in_R3_C1_dqdPE2 = minv[2][0];
        minv_block_in_R4_C1_dqdPE2 = minv[3][0];
        minv_block_in_R5_C1_dqdPE2 = minv[4][0];
        minv_block_in_R6_C1_dqdPE2 = minv[5][0];
        minv_block_in_R7_C1_dqdPE2 = minv[6][0];

        minv_block_in_R1_C2_dqdPE2 = minv[0][1];
        minv_block_in_R2_C2_dqdPE2 = minv[1][1];
        minv_block_in_R3_C2_dqdPE2 = minv[2][1];
        minv_block_in_R4_C2_dqdPE2 = minv[3][1];
        minv_block_in_R5_C2_dqdPE2 = minv[4][1];
        minv_block_in_R6_C2_dqdPE2 = minv[5][1];
        minv_block_in_R7_C2_dqdPE2 = minv[6][1];

        minv_block_in_R1_C3_dqdPE2 = minv[0][2];
        minv_block_in_R2_C3_dqdPE2 = minv[1][2];
        minv_block_in_R3_C3_dqdPE2 = minv[2][2];
        minv_block_in_R4_C3_dqdPE2 = minv[3][2];
        minv_block_in_R5_C3_dqdPE2 = minv[4][2];
        minv_block_in_R6_C3_dqdPE2 = minv[5][2];
        minv_block_in_R7_C3_dqdPE2 = minv[6][2];

        minv_block_in_R1_C4_dqdPE2 = minv[0][3];
        minv_block_in_R2_C4_dqdPE2 = minv[1][3];
        minv_block_in_R3_C4_dqdPE2 = minv[2][3];
        minv_block_in_R4_C4_dqdPE2 = minv[3][3];
        minv_block_in_R5_C4_dqdPE2 = minv[4][3];
        minv_block_in_R6_C4_dqdPE2 = minv[5][3];
        minv_block_in_R7_C4_dqdPE2 = minv[6][3];

        minv_block_in_R1_C5_dqdPE2 = minv[0][4];
        minv_block_in_R2_C5_dqdPE2 = minv[1][4];
        minv_block_in_R3_C5_dqdPE2 = minv[2][4];
        minv_block_in_R4_C5_dqdPE2 = minv[3][4];
        minv_block_in_R5_C5_dqdPE2 = minv[4][4];
        minv_block_in_R6_C5_dqdPE2 = minv[5][4];
        minv_block_in_R7_C5_dqdPE2 = minv[6][4];

        minv_block_in_R1_C6_dqdPE2 = minv[0][5];
        minv_block_in_R2_C6_dqdPE2 = minv[1][5];
        minv_block_in_R3_C6_dqdPE2 = minv[2][5];
        minv_block_in_R4_C6_dqdPE2 = minv[3][5];
        minv_block_in_R5_C6_dqdPE2 = minv[4][5];
        minv_block_in_R6_C6_dqdPE2 = minv[5][5];
        minv_block_in_R7_C6_dqdPE2 = minv[6][5];

        minv_block_in_R1_C7_dqdPE2 = minv[0][6];
        minv_block_in_R2_C7_dqdPE2 = minv[1][6];
        minv_block_in_R3_C7_dqdPE2 = minv[2][6];
        minv_block_in_R4_C7_dqdPE2 = minv[3][6];
        minv_block_in_R5_C7_dqdPE2 = minv[4][6];
        minv_block_in_R6_C7_dqdPE2 = minv[5][6];
        minv_block_in_R7_C7_dqdPE2 = minv[6][6];

        minv_block_in_R1_C1_dqdPE3 = minv[0][0];
        minv_block_in_R2_C1_dqdPE3 = minv[1][0];
        minv_block_in_R3_C1_dqdPE3 = minv[2][0];
        minv_block_in_R4_C1_dqdPE3 = minv[3][0];
        minv_block_in_R5_C1_dqdPE3 = minv[4][0];
        minv_block_in_R6_C1_dqdPE3 = minv[5][0];
        minv_block_in_R7_C1_dqdPE3 = minv[6][0];

        minv_block_in_R1_C2_dqdPE3 = minv[0][1];
        minv_block_in_R2_C2_dqdPE3 = minv[1][1];
        minv_block_in_R3_C2_dqdPE3 = minv[2][1];
        minv_block_in_R4_C2_dqdPE3 = minv[3][1];
        minv_block_in_R5_C2_dqdPE3 = minv[4][1];
        minv_block_in_R6_C2_dqdPE3 = minv[5][1];
        minv_block_in_R7_C2_dqdPE3 = minv[6][1];

        minv_block_in_R1_C3_dqdPE3 = minv[0][2];
        minv_block_in_R2_C3_dqdPE3 = minv[1][2];
        minv_block_in_R3_C3_dqdPE3 = minv[2][2];
        minv_block_in_R4_C3_dqdPE3 = minv[3][2];
        minv_block_in_R5_C3_dqdPE3 = minv[4][2];
        minv_block_in_R6_C3_dqdPE3 = minv[5][2];
        minv_block_in_R7_C3_dqdPE3 = minv[6][2];

        minv_block_in_R1_C4_dqdPE3 = minv[0][3];
        minv_block_in_R2_C4_dqdPE3 = minv[1][3];
        minv_block_in_R3_C4_dqdPE3 = minv[2][3];
        minv_block_in_R4_C4_dqdPE3 = minv[3][3];
        minv_block_in_R5_C4_dqdPE3 = minv[4][3];
        minv_block_in_R6_C4_dqdPE3 = minv[5][3];
        minv_block_in_R7_C4_dqdPE3 = minv[6][3];

        minv_block_in_R1_C5_dqdPE3 = minv[0][4];
        minv_block_in_R2_C5_dqdPE3 = minv[1][4];
        minv_block_in_R3_C5_dqdPE3 = minv[2][4];
        minv_block_in_R4_C5_dqdPE3 = minv[3][4];
        minv_block_in_R5_C5_dqdPE3 = minv[4][4];
        minv_block_in_R6_C5_dqdPE3 = minv[5][4];
        minv_block_in_R7_C5_dqdPE3 = minv[6][4];

        minv_block_in_R1_C6_dqdPE3 = minv[0][5];
        minv_block_in_R2_C6_dqdPE3 = minv[1][5];
        minv_block_in_R3_C6_dqdPE3 = minv[2][5];
        minv_block_in_R4_C6_dqdPE3 = minv[3][5];
        minv_block_in_R5_C6_dqdPE3 = minv[4][5];
        minv_block_in_R6_C6_dqdPE3 = minv[5][5];
        minv_block_in_R7_C6_dqdPE3 = minv[6][5];

        minv_block_in_R1_C7_dqdPE3 = minv[0][6];
        minv_block_in_R2_C7_dqdPE3 = minv[1][6];
        minv_block_in_R3_C7_dqdPE3 = minv[2][6];
        minv_block_in_R4_C7_dqdPE3 = minv[3][6];
        minv_block_in_R5_C7_dqdPE3 = minv[4][6];
        minv_block_in_R6_C7_dqdPE3 = minv[5][6];
        minv_block_in_R7_C7_dqdPE3 = minv[6][6];

        minv_block_in_R1_C1_dqdPE4 = minv[0][0];
        minv_block_in_R2_C1_dqdPE4 = minv[1][0];
        minv_block_in_R3_C1_dqdPE4 = minv[2][0];
        minv_block_in_R4_C1_dqdPE4 = minv[3][0];
        minv_block_in_R5_C1_dqdPE4 = minv[4][0];
        minv_block_in_R6_C1_dqdPE4 = minv[5][0];
        minv_block_in_R7_C1_dqdPE4 = minv[6][0];

        minv_block_in_R1_C2_dqdPE4 = minv[0][1];
        minv_block_in_R2_C2_dqdPE4 = minv[1][1];
        minv_block_in_R3_C2_dqdPE4 = minv[2][1];
        minv_block_in_R4_C2_dqdPE4 = minv[3][1];
        minv_block_in_R5_C2_dqdPE4 = minv[4][1];
        minv_block_in_R6_C2_dqdPE4 = minv[5][1];
        minv_block_in_R7_C2_dqdPE4 = minv[6][1];

        minv_block_in_R1_C3_dqdPE4 = minv[0][2];
        minv_block_in_R2_C3_dqdPE4 = minv[1][2];
        minv_block_in_R3_C3_dqdPE4 = minv[2][2];
        minv_block_in_R4_C3_dqdPE4 = minv[3][2];
        minv_block_in_R5_C3_dqdPE4 = minv[4][2];
        minv_block_in_R6_C3_dqdPE4 = minv[5][2];
        minv_block_in_R7_C3_dqdPE4 = minv[6][2];

        minv_block_in_R1_C4_dqdPE4 = minv[0][3];
        minv_block_in_R2_C4_dqdPE4 = minv[1][3];
        minv_block_in_R3_C4_dqdPE4 = minv[2][3];
        minv_block_in_R4_C4_dqdPE4 = minv[3][3];
        minv_block_in_R5_C4_dqdPE4 = minv[4][3];
        minv_block_in_R6_C4_dqdPE4 = minv[5][3];
        minv_block_in_R7_C4_dqdPE4 = minv[6][3];

        minv_block_in_R1_C5_dqdPE4 = minv[0][4];
        minv_block_in_R2_C5_dqdPE4 = minv[1][4];
        minv_block_in_R3_C5_dqdPE4 = minv[2][4];
        minv_block_in_R4_C5_dqdPE4 = minv[3][4];
        minv_block_in_R5_C5_dqdPE4 = minv[4][4];
        minv_block_in_R6_C5_dqdPE4 = minv[5][4];
        minv_block_in_R7_C5_dqdPE4 = minv[6][4];

        minv_block_in_R1_C6_dqdPE4 = minv[0][5];
        minv_block_in_R2_C6_dqdPE4 = minv[1][5];
        minv_block_in_R3_C6_dqdPE4 = minv[2][5];
        minv_block_in_R4_C6_dqdPE4 = minv[3][5];
        minv_block_in_R5_C6_dqdPE4 = minv[4][5];
        minv_block_in_R6_C6_dqdPE4 = minv[5][5];
        minv_block_in_R7_C6_dqdPE4 = minv[6][5];

        minv_block_in_R1_C7_dqdPE4 = minv[0][6];
        minv_block_in_R2_C7_dqdPE4 = minv[1][6];
        minv_block_in_R3_C7_dqdPE4 = minv[2][6];
        minv_block_in_R4_C7_dqdPE4 = minv[3][6];
        minv_block_in_R5_C7_dqdPE4 = minv[4][6];
        minv_block_in_R6_C7_dqdPE4 = minv[5][6];
        minv_block_in_R7_C7_dqdPE4 = minv[6][6];

        minv_block_in_R1_C1_dqdPE5 = minv[0][0];
        minv_block_in_R2_C1_dqdPE5 = minv[1][0];
        minv_block_in_R3_C1_dqdPE5 = minv[2][0];
        minv_block_in_R4_C1_dqdPE5 = minv[3][0];
        minv_block_in_R5_C1_dqdPE5 = minv[4][0];
        minv_block_in_R6_C1_dqdPE5 = minv[5][0];
        minv_block_in_R7_C1_dqdPE5 = minv[6][0];

        minv_block_in_R1_C2_dqdPE5 = minv[0][1];
        minv_block_in_R2_C2_dqdPE5 = minv[1][1];
        minv_block_in_R3_C2_dqdPE5 = minv[2][1];
        minv_block_in_R4_C2_dqdPE5 = minv[3][1];
        minv_block_in_R5_C2_dqdPE5 = minv[4][1];
        minv_block_in_R6_C2_dqdPE5 = minv[5][1];
        minv_block_in_R7_C2_dqdPE5 = minv[6][1];

        minv_block_in_R1_C3_dqdPE5 = minv[0][2];
        minv_block_in_R2_C3_dqdPE5 = minv[1][2];
        minv_block_in_R3_C3_dqdPE5 = minv[2][2];
        minv_block_in_R4_C3_dqdPE5 = minv[3][2];
        minv_block_in_R5_C3_dqdPE5 = minv[4][2];
        minv_block_in_R6_C3_dqdPE5 = minv[5][2];
        minv_block_in_R7_C3_dqdPE5 = minv[6][2];

        minv_block_in_R1_C4_dqdPE5 = minv[0][3];
        minv_block_in_R2_C4_dqdPE5 = minv[1][3];
        minv_block_in_R3_C4_dqdPE5 = minv[2][3];
        minv_block_in_R4_C4_dqdPE5 = minv[3][3];
        minv_block_in_R5_C4_dqdPE5 = minv[4][3];
        minv_block_in_R6_C4_dqdPE5 = minv[5][3];
        minv_block_in_R7_C4_dqdPE5 = minv[6][3];

        minv_block_in_R1_C5_dqdPE5 = minv[0][4];
        minv_block_in_R2_C5_dqdPE5 = minv[1][4];
        minv_block_in_R3_C5_dqdPE5 = minv[2][4];
        minv_block_in_R4_C5_dqdPE5 = minv[3][4];
        minv_block_in_R5_C5_dqdPE5 = minv[4][4];
        minv_block_in_R6_C5_dqdPE5 = minv[5][4];
        minv_block_in_R7_C5_dqdPE5 = minv[6][4];

        minv_block_in_R1_C6_dqdPE5 = minv[0][5];
        minv_block_in_R2_C6_dqdPE5 = minv[1][5];
        minv_block_in_R3_C6_dqdPE5 = minv[2][5];
        minv_block_in_R4_C6_dqdPE5 = minv[3][5];
        minv_block_in_R5_C6_dqdPE5 = minv[4][5];
        minv_block_in_R6_C6_dqdPE5 = minv[5][5];
        minv_block_in_R7_C6_dqdPE5 = minv[6][5];

        minv_block_in_R1_C7_dqdPE5 = minv[0][6];
        minv_block_in_R2_C7_dqdPE5 = minv[1][6];
        minv_block_in_R3_C7_dqdPE5 = minv[2][6];
        minv_block_in_R4_C7_dqdPE5 = minv[3][6];
        minv_block_in_R5_C7_dqdPE5 = minv[4][6];
        minv_block_in_R6_C7_dqdPE5 = minv[5][6];
        minv_block_in_R7_C7_dqdPE5 = minv[6][6];

        minv_block_in_R1_C1_dqdPE6 = minv[0][0];
        minv_block_in_R2_C1_dqdPE6 = minv[1][0];
        minv_block_in_R3_C1_dqdPE6 = minv[2][0];
        minv_block_in_R4_C1_dqdPE6 = minv[3][0];
        minv_block_in_R5_C1_dqdPE6 = minv[4][0];
        minv_block_in_R6_C1_dqdPE6 = minv[5][0];
        minv_block_in_R7_C1_dqdPE6 = minv[6][0];

        minv_block_in_R1_C2_dqdPE6 = minv[0][1];
        minv_block_in_R2_C2_dqdPE6 = minv[1][1];
        minv_block_in_R3_C2_dqdPE6 = minv[2][1];
        minv_block_in_R4_C2_dqdPE6 = minv[3][1];
        minv_block_in_R5_C2_dqdPE6 = minv[4][1];
        minv_block_in_R6_C2_dqdPE6 = minv[5][1];
        minv_block_in_R7_C2_dqdPE6 = minv[6][1];

        minv_block_in_R1_C3_dqdPE6 = minv[0][2];
        minv_block_in_R2_C3_dqdPE6 = minv[1][2];
        minv_block_in_R3_C3_dqdPE6 = minv[2][2];
        minv_block_in_R4_C3_dqdPE6 = minv[3][2];
        minv_block_in_R5_C3_dqdPE6 = minv[4][2];
        minv_block_in_R6_C3_dqdPE6 = minv[5][2];
        minv_block_in_R7_C3_dqdPE6 = minv[6][2];

        minv_block_in_R1_C4_dqdPE6 = minv[0][3];
        minv_block_in_R2_C4_dqdPE6 = minv[1][3];
        minv_block_in_R3_C4_dqdPE6 = minv[2][3];
        minv_block_in_R4_C4_dqdPE6 = minv[3][3];
        minv_block_in_R5_C4_dqdPE6 = minv[4][3];
        minv_block_in_R6_C4_dqdPE6 = minv[5][3];
        minv_block_in_R7_C4_dqdPE6 = minv[6][3];

        minv_block_in_R1_C5_dqdPE6 = minv[0][4];
        minv_block_in_R2_C5_dqdPE6 = minv[1][4];
        minv_block_in_R3_C5_dqdPE6 = minv[2][4];
        minv_block_in_R4_C5_dqdPE6 = minv[3][4];
        minv_block_in_R5_C5_dqdPE6 = minv[4][4];
        minv_block_in_R6_C5_dqdPE6 = minv[5][4];
        minv_block_in_R7_C5_dqdPE6 = minv[6][4];

        minv_block_in_R1_C6_dqdPE6 = minv[0][5];
        minv_block_in_R2_C6_dqdPE6 = minv[1][5];
        minv_block_in_R3_C6_dqdPE6 = minv[2][5];
        minv_block_in_R4_C6_dqdPE6 = minv[3][5];
        minv_block_in_R5_C6_dqdPE6 = minv[4][5];
        minv_block_in_R6_C6_dqdPE6 = minv[5][5];
        minv_block_in_R7_C6_dqdPE6 = minv[6][5];

        minv_block_in_R1_C7_dqdPE6 = minv[0][6];
        minv_block_in_R2_C7_dqdPE6 = minv[1][6];
        minv_block_in_R3_C7_dqdPE6 = minv[2][6];
        minv_block_in_R4_C7_dqdPE6 = minv[3][6];
        minv_block_in_R5_C7_dqdPE6 = minv[4][6];
        minv_block_in_R6_C7_dqdPE6 = minv[5][6];
        minv_block_in_R7_C7_dqdPE6 = minv[6][6];

        minv_block_in_R1_C1_dqdPE7 = minv[0][0];
        minv_block_in_R2_C1_dqdPE7 = minv[1][0];
        minv_block_in_R3_C1_dqdPE7 = minv[2][0];
        minv_block_in_R4_C1_dqdPE7 = minv[3][0];
        minv_block_in_R5_C1_dqdPE7 = minv[4][0];
        minv_block_in_R6_C1_dqdPE7 = minv[5][0];
        minv_block_in_R7_C1_dqdPE7 = minv[6][0];

        minv_block_in_R1_C2_dqdPE7 = minv[0][1];
        minv_block_in_R2_C2_dqdPE7 = minv[1][1];
        minv_block_in_R3_C2_dqdPE7 = minv[2][1];
        minv_block_in_R4_C2_dqdPE7 = minv[3][1];
        minv_block_in_R5_C2_dqdPE7 = minv[4][1];
        minv_block_in_R6_C2_dqdPE7 = minv[5][1];
        minv_block_in_R7_C2_dqdPE7 = minv[6][1];

        minv_block_in_R1_C3_dqdPE7 = minv[0][2];
        minv_block_in_R2_C3_dqdPE7 = minv[1][2];
        minv_block_in_R3_C3_dqdPE7 = minv[2][2];
        minv_block_in_R4_C3_dqdPE7 = minv[3][2];
        minv_block_in_R5_C3_dqdPE7 = minv[4][2];
        minv_block_in_R6_C3_dqdPE7 = minv[5][2];
        minv_block_in_R7_C3_dqdPE7 = minv[6][2];

        minv_block_in_R1_C4_dqdPE7 = minv[0][3];
        minv_block_in_R2_C4_dqdPE7 = minv[1][3];
        minv_block_in_R3_C4_dqdPE7 = minv[2][3];
        minv_block_in_R4_C4_dqdPE7 = minv[3][3];
        minv_block_in_R5_C4_dqdPE7 = minv[4][3];
        minv_block_in_R6_C4_dqdPE7 = minv[5][3];
        minv_block_in_R7_C4_dqdPE7 = minv[6][3];

        minv_block_in_R1_C5_dqdPE7 = minv[0][4];
        minv_block_in_R2_C5_dqdPE7 = minv[1][4];
        minv_block_in_R3_C5_dqdPE7 = minv[2][4];
        minv_block_in_R4_C5_dqdPE7 = minv[3][4];
        minv_block_in_R5_C5_dqdPE7 = minv[4][4];
        minv_block_in_R6_C5_dqdPE7 = minv[5][4];
        minv_block_in_R7_C5_dqdPE7 = minv[6][4];

        minv_block_in_R1_C6_dqdPE7 = minv[0][5];
        minv_block_in_R2_C6_dqdPE7 = minv[1][5];
        minv_block_in_R3_C6_dqdPE7 = minv[2][5];
        minv_block_in_R4_C6_dqdPE7 = minv[3][5];
        minv_block_in_R5_C6_dqdPE7 = minv[4][5];
        minv_block_in_R6_C6_dqdPE7 = minv[5][5];
        minv_block_in_R7_C6_dqdPE7 = minv[6][5];

        minv_block_in_R1_C7_dqdPE7 = minv[0][6];
        minv_block_in_R2_C7_dqdPE7 = minv[1][6];
        minv_block_in_R3_C7_dqdPE7 = minv[2][6];
        minv_block_in_R4_C7_dqdPE7 = minv[3][6];
        minv_block_in_R5_C7_dqdPE7 = minv[4][6];
        minv_block_in_R6_C7_dqdPE7 = minv[5][6];
        minv_block_in_R7_C7_dqdPE7 = minv[6][6];

        dtau_vec_in_R1_dqdPE1 = dtau_mat_curr[0][0];
        dtau_vec_in_R2_dqdPE1 = dtau_mat_curr[1][0];
        dtau_vec_in_R3_dqdPE1 = dtau_mat_curr[2][0];
        dtau_vec_in_R4_dqdPE1 = dtau_mat_curr[3][0];
        dtau_vec_in_R5_dqdPE1 = dtau_mat_curr[4][0];
        dtau_vec_in_R6_dqdPE1 = dtau_mat_curr[5][0];
        dtau_vec_in_R7_dqdPE1 = dtau_mat_curr[6][0];

        dtau_vec_in_R1_dqdPE2 = dtau_mat_curr[0][1];
        dtau_vec_in_R2_dqdPE2 = dtau_mat_curr[1][1];
        dtau_vec_in_R3_dqdPE2 = dtau_mat_curr[2][1];
        dtau_vec_in_R4_dqdPE2 = dtau_mat_curr[3][1];
        dtau_vec_in_R5_dqdPE2 = dtau_mat_curr[4][1];
        dtau_vec_in_R6_dqdPE2 = dtau_mat_curr[5][1];
        dtau_vec_in_R7_dqdPE2 = dtau_mat_curr[6][1];

        dtau_vec_in_R1_dqdPE3 = dtau_mat_curr[0][2];
        dtau_vec_in_R2_dqdPE3 = dtau_mat_curr[1][2];
        dtau_vec_in_R3_dqdPE3 = dtau_mat_curr[2][2];
        dtau_vec_in_R4_dqdPE3 = dtau_mat_curr[3][2];
        dtau_vec_in_R5_dqdPE3 = dtau_mat_curr[4][2];
        dtau_vec_in_R6_dqdPE3 = dtau_mat_curr[5][2];
        dtau_vec_in_R7_dqdPE3 = dtau_mat_curr[6][2];

        dtau_vec_in_R1_dqdPE4 = dtau_mat_curr[0][3];
        dtau_vec_in_R2_dqdPE4 = dtau_mat_curr[1][3];
        dtau_vec_in_R3_dqdPE4 = dtau_mat_curr[2][3];
        dtau_vec_in_R4_dqdPE4 = dtau_mat_curr[3][3];
        dtau_vec_in_R5_dqdPE4 = dtau_mat_curr[4][3];
        dtau_vec_in_R6_dqdPE4 = dtau_mat_curr[5][3];
        dtau_vec_in_R7_dqdPE4 = dtau_mat_curr[6][3];

        dtau_vec_in_R1_dqdPE5 = dtau_mat_curr[0][4];
        dtau_vec_in_R2_dqdPE5 = dtau_mat_curr[1][4];
        dtau_vec_in_R3_dqdPE5 = dtau_mat_curr[2][4];
        dtau_vec_in_R4_dqdPE5 = dtau_mat_curr[3][4];
        dtau_vec_in_R5_dqdPE5 = dtau_mat_curr[4][4];
        dtau_vec_in_R6_dqdPE5 = dtau_mat_curr[5][4];
        dtau_vec_in_R7_dqdPE5 = dtau_mat_curr[6][4];

        dtau_vec_in_R1_dqdPE6 = dtau_mat_curr[0][5];
        dtau_vec_in_R2_dqdPE6 = dtau_mat_curr[1][5];
        dtau_vec_in_R3_dqdPE6 = dtau_mat_curr[2][5];
        dtau_vec_in_R4_dqdPE6 = dtau_mat_curr[3][5];
        dtau_vec_in_R5_dqdPE6 = dtau_mat_curr[4][5];
        dtau_vec_in_R6_dqdPE6 = dtau_mat_curr[5][5];
        dtau_vec_in_R7_dqdPE6 = dtau_mat_curr[6][5];

        dtau_vec_in_R1_dqdPE7 = dtau_mat_curr[0][6];
        dtau_vec_in_R2_dqdPE7 = dtau_mat_curr[1][6];
        dtau_vec_in_R3_dqdPE7 = dtau_mat_curr[2][6];
        dtau_vec_in_R4_dqdPE7 = dtau_mat_curr[3][6];
        dtau_vec_in_R5_dqdPE7 = dtau_mat_curr[4][6];
        dtau_vec_in_R6_dqdPE7 = dtau_mat_curr[5][6];
        dtau_vec_in_R7_dqdPE7 = dtau_mat_curr[6][6];

    end

endcase

bproc.minv_block_in_R1_C1_dqdPE1(minv_block_in_R1_C1_dqdPE1);
bproc.minv_block_in_R2_C1_dqdPE1(minv_block_in_R2_C1_dqdPE1);
bproc.minv_block_in_R3_C1_dqdPE1(minv_block_in_R3_C1_dqdPE1);
bproc.minv_block_in_R4_C1_dqdPE1(minv_block_in_R4_C1_dqdPE1);
bproc.minv_block_in_R5_C1_dqdPE1(minv_block_in_R5_C1_dqdPE1);
bproc.minv_block_in_R6_C1_dqdPE1(minv_block_in_R6_C1_dqdPE1);
bproc.minv_block_in_R7_C1_dqdPE1(minv_block_in_R7_C1_dqdPE1);

bproc.minv_block_in_R1_C2_dqdPE1(minv_block_in_R1_C2_dqdPE1);
bproc.minv_block_in_R2_C2_dqdPE1(minv_block_in_R2_C2_dqdPE1);
bproc.minv_block_in_R3_C2_dqdPE1(minv_block_in_R3_C2_dqdPE1);
bproc.minv_block_in_R4_C2_dqdPE1(minv_block_in_R4_C2_dqdPE1);
bproc.minv_block_in_R5_C2_dqdPE1(minv_block_in_R5_C2_dqdPE1);
bproc.minv_block_in_R6_C2_dqdPE1(minv_block_in_R6_C2_dqdPE1);
bproc.minv_block_in_R7_C2_dqdPE1(minv_block_in_R7_C2_dqdPE1);

bproc.minv_block_in_R1_C3_dqdPE1(minv_block_in_R1_C3_dqdPE1);
bproc.minv_block_in_R2_C3_dqdPE1(minv_block_in_R2_C3_dqdPE1);
bproc.minv_block_in_R3_C3_dqdPE1(minv_block_in_R3_C3_dqdPE1);
bproc.minv_block_in_R4_C3_dqdPE1(minv_block_in_R4_C3_dqdPE1);
bproc.minv_block_in_R5_C3_dqdPE1(minv_block_in_R5_C3_dqdPE1);
bproc.minv_block_in_R6_C3_dqdPE1(minv_block_in_R6_C3_dqdPE1);
bproc.minv_block_in_R7_C3_dqdPE1(minv_block_in_R7_C3_dqdPE1);

bproc.minv_block_in_R1_C4_dqdPE1(minv_block_in_R1_C4_dqdPE1);
bproc.minv_block_in_R2_C4_dqdPE1(minv_block_in_R2_C4_dqdPE1);
bproc.minv_block_in_R3_C4_dqdPE1(minv_block_in_R3_C4_dqdPE1);
bproc.minv_block_in_R4_C4_dqdPE1(minv_block_in_R4_C4_dqdPE1);
bproc.minv_block_in_R5_C4_dqdPE1(minv_block_in_R5_C4_dqdPE1);
bproc.minv_block_in_R6_C4_dqdPE1(minv_block_in_R6_C4_dqdPE1);
bproc.minv_block_in_R7_C4_dqdPE1(minv_block_in_R7_C4_dqdPE1);

bproc.minv_block_in_R1_C5_dqdPE1(minv_block_in_R1_C5_dqdPE1);
bproc.minv_block_in_R2_C5_dqdPE1(minv_block_in_R2_C5_dqdPE1);
bproc.minv_block_in_R3_C5_dqdPE1(minv_block_in_R3_C5_dqdPE1);
bproc.minv_block_in_R4_C5_dqdPE1(minv_block_in_R4_C5_dqdPE1);
bproc.minv_block_in_R5_C5_dqdPE1(minv_block_in_R5_C5_dqdPE1);
bproc.minv_block_in_R6_C5_dqdPE1(minv_block_in_R6_C5_dqdPE1);
bproc.minv_block_in_R7_C5_dqdPE1(minv_block_in_R7_C5_dqdPE1);

bproc.minv_block_in_R1_C6_dqdPE1(minv_block_in_R1_C6_dqdPE1);
bproc.minv_block_in_R2_C6_dqdPE1(minv_block_in_R2_C6_dqdPE1);
bproc.minv_block_in_R3_C6_dqdPE1(minv_block_in_R3_C6_dqdPE1);
bproc.minv_block_in_R4_C6_dqdPE1(minv_block_in_R4_C6_dqdPE1);
bproc.minv_block_in_R5_C6_dqdPE1(minv_block_in_R5_C6_dqdPE1);
bproc.minv_block_in_R6_C6_dqdPE1(minv_block_in_R6_C6_dqdPE1);
bproc.minv_block_in_R7_C6_dqdPE1(minv_block_in_R7_C6_dqdPE1);

bproc.minv_block_in_R1_C7_dqdPE1(minv_block_in_R1_C7_dqdPE1);
bproc.minv_block_in_R2_C7_dqdPE1(minv_block_in_R2_C7_dqdPE1);
bproc.minv_block_in_R3_C7_dqdPE1(minv_block_in_R3_C7_dqdPE1);
bproc.minv_block_in_R4_C7_dqdPE1(minv_block_in_R4_C7_dqdPE1);
bproc.minv_block_in_R5_C7_dqdPE1(minv_block_in_R5_C7_dqdPE1);
bproc.minv_block_in_R6_C7_dqdPE1(minv_block_in_R6_C7_dqdPE1);
bproc.minv_block_in_R7_C7_dqdPE1(minv_block_in_R7_C7_dqdPE1);

bproc.dtau_vec_in_R1_dqdPE1(dtau_vec_in_R1_dqdPE1);
bproc.dtau_vec_in_R2_dqdPE1(dtau_vec_in_R2_dqdPE1);
bproc.dtau_vec_in_R3_dqdPE1(dtau_vec_in_R3_dqdPE1);
bproc.dtau_vec_in_R4_dqdPE1(dtau_vec_in_R4_dqdPE1);
bproc.dtau_vec_in_R5_dqdPE1(dtau_vec_in_R5_dqdPE1);
bproc.dtau_vec_in_R6_dqdPE1(dtau_vec_in_R6_dqdPE1);
bproc.dtau_vec_in_R7_dqdPE1(dtau_vec_in_R7_dqdPE1);

bproc.minv_block_in_R1_C1_dqdPE2(minv_block_in_R1_C1_dqdPE2);
bproc.minv_block_in_R2_C1_dqdPE2(minv_block_in_R2_C1_dqdPE2);
bproc.minv_block_in_R3_C1_dqdPE2(minv_block_in_R3_C1_dqdPE2);
bproc.minv_block_in_R4_C1_dqdPE2(minv_block_in_R4_C1_dqdPE2);
bproc.minv_block_in_R5_C1_dqdPE2(minv_block_in_R5_C1_dqdPE2);
bproc.minv_block_in_R6_C1_dqdPE2(minv_block_in_R6_C1_dqdPE2);
bproc.minv_block_in_R7_C1_dqdPE2(minv_block_in_R7_C1_dqdPE2);

bproc.minv_block_in_R1_C2_dqdPE2(minv_block_in_R1_C2_dqdPE2);
bproc.minv_block_in_R2_C2_dqdPE2(minv_block_in_R2_C2_dqdPE2);
bproc.minv_block_in_R3_C2_dqdPE2(minv_block_in_R3_C2_dqdPE2);
bproc.minv_block_in_R4_C2_dqdPE2(minv_block_in_R4_C2_dqdPE2);
bproc.minv_block_in_R5_C2_dqdPE2(minv_block_in_R5_C2_dqdPE2);
bproc.minv_block_in_R6_C2_dqdPE2(minv_block_in_R6_C2_dqdPE2);
bproc.minv_block_in_R7_C2_dqdPE2(minv_block_in_R7_C2_dqdPE2);

bproc.minv_block_in_R1_C3_dqdPE2(minv_block_in_R1_C3_dqdPE2);
bproc.minv_block_in_R2_C3_dqdPE2(minv_block_in_R2_C3_dqdPE2);
bproc.minv_block_in_R3_C3_dqdPE2(minv_block_in_R3_C3_dqdPE2);
bproc.minv_block_in_R4_C3_dqdPE2(minv_block_in_R4_C3_dqdPE2);
bproc.minv_block_in_R5_C3_dqdPE2(minv_block_in_R5_C3_dqdPE2);
bproc.minv_block_in_R6_C3_dqdPE2(minv_block_in_R6_C3_dqdPE2);
bproc.minv_block_in_R7_C3_dqdPE2(minv_block_in_R7_C3_dqdPE2);

bproc.minv_block_in_R1_C4_dqdPE2(minv_block_in_R1_C4_dqdPE2);
bproc.minv_block_in_R2_C4_dqdPE2(minv_block_in_R2_C4_dqdPE2);
bproc.minv_block_in_R3_C4_dqdPE2(minv_block_in_R3_C4_dqdPE2);
bproc.minv_block_in_R4_C4_dqdPE2(minv_block_in_R4_C4_dqdPE2);
bproc.minv_block_in_R5_C4_dqdPE2(minv_block_in_R5_C4_dqdPE2);
bproc.minv_block_in_R6_C4_dqdPE2(minv_block_in_R6_C4_dqdPE2);
bproc.minv_block_in_R7_C4_dqdPE2(minv_block_in_R7_C4_dqdPE2);

bproc.minv_block_in_R1_C5_dqdPE2(minv_block_in_R1_C5_dqdPE2);
bproc.minv_block_in_R2_C5_dqdPE2(minv_block_in_R2_C5_dqdPE2);
bproc.minv_block_in_R3_C5_dqdPE2(minv_block_in_R3_C5_dqdPE2);
bproc.minv_block_in_R4_C5_dqdPE2(minv_block_in_R4_C5_dqdPE2);
bproc.minv_block_in_R5_C5_dqdPE2(minv_block_in_R5_C5_dqdPE2);
bproc.minv_block_in_R6_C5_dqdPE2(minv_block_in_R6_C5_dqdPE2);
bproc.minv_block_in_R7_C5_dqdPE2(minv_block_in_R7_C5_dqdPE2);

bproc.minv_block_in_R1_C6_dqdPE2(minv_block_in_R1_C6_dqdPE2);
bproc.minv_block_in_R2_C6_dqdPE2(minv_block_in_R2_C6_dqdPE2);
bproc.minv_block_in_R3_C6_dqdPE2(minv_block_in_R3_C6_dqdPE2);
bproc.minv_block_in_R4_C6_dqdPE2(minv_block_in_R4_C6_dqdPE2);
bproc.minv_block_in_R5_C6_dqdPE2(minv_block_in_R5_C6_dqdPE2);
bproc.minv_block_in_R6_C6_dqdPE2(minv_block_in_R6_C6_dqdPE2);
bproc.minv_block_in_R7_C6_dqdPE2(minv_block_in_R7_C6_dqdPE2);

bproc.minv_block_in_R1_C7_dqdPE2(minv_block_in_R1_C7_dqdPE2);
bproc.minv_block_in_R2_C7_dqdPE2(minv_block_in_R2_C7_dqdPE2);
bproc.minv_block_in_R3_C7_dqdPE2(minv_block_in_R3_C7_dqdPE2);
bproc.minv_block_in_R4_C7_dqdPE2(minv_block_in_R4_C7_dqdPE2);
bproc.minv_block_in_R5_C7_dqdPE2(minv_block_in_R5_C7_dqdPE2);
bproc.minv_block_in_R6_C7_dqdPE2(minv_block_in_R6_C7_dqdPE2);
bproc.minv_block_in_R7_C7_dqdPE2(minv_block_in_R7_C7_dqdPE2);

bproc.dtau_vec_in_R1_dqdPE2(dtau_vec_in_R1_dqdPE2);
bproc.dtau_vec_in_R2_dqdPE2(dtau_vec_in_R2_dqdPE2);
bproc.dtau_vec_in_R3_dqdPE2(dtau_vec_in_R3_dqdPE2);
bproc.dtau_vec_in_R4_dqdPE2(dtau_vec_in_R4_dqdPE2);
bproc.dtau_vec_in_R5_dqdPE2(dtau_vec_in_R5_dqdPE2);
bproc.dtau_vec_in_R6_dqdPE2(dtau_vec_in_R6_dqdPE2);
bproc.dtau_vec_in_R7_dqdPE2(dtau_vec_in_R7_dqdPE2);

bproc.minv_block_in_R1_C1_dqdPE3(minv_block_in_R1_C1_dqdPE3);
bproc.minv_block_in_R2_C1_dqdPE3(minv_block_in_R2_C1_dqdPE3);
bproc.minv_block_in_R3_C1_dqdPE3(minv_block_in_R3_C1_dqdPE3);
bproc.minv_block_in_R4_C1_dqdPE3(minv_block_in_R4_C1_dqdPE3);
bproc.minv_block_in_R5_C1_dqdPE3(minv_block_in_R5_C1_dqdPE3);
bproc.minv_block_in_R6_C1_dqdPE3(minv_block_in_R6_C1_dqdPE3);
bproc.minv_block_in_R7_C1_dqdPE3(minv_block_in_R7_C1_dqdPE3);

bproc.minv_block_in_R1_C2_dqdPE3(minv_block_in_R1_C2_dqdPE3);
bproc.minv_block_in_R2_C2_dqdPE3(minv_block_in_R2_C2_dqdPE3);
bproc.minv_block_in_R3_C2_dqdPE3(minv_block_in_R3_C2_dqdPE3);
bproc.minv_block_in_R4_C2_dqdPE3(minv_block_in_R4_C2_dqdPE3);
bproc.minv_block_in_R5_C2_dqdPE3(minv_block_in_R5_C2_dqdPE3);
bproc.minv_block_in_R6_C2_dqdPE3(minv_block_in_R6_C2_dqdPE3);
bproc.minv_block_in_R7_C2_dqdPE3(minv_block_in_R7_C2_dqdPE3);

bproc.minv_block_in_R1_C3_dqdPE3(minv_block_in_R1_C3_dqdPE3);
bproc.minv_block_in_R2_C3_dqdPE3(minv_block_in_R2_C3_dqdPE3);
bproc.minv_block_in_R3_C3_dqdPE3(minv_block_in_R3_C3_dqdPE3);
bproc.minv_block_in_R4_C3_dqdPE3(minv_block_in_R4_C3_dqdPE3);
bproc.minv_block_in_R5_C3_dqdPE3(minv_block_in_R5_C3_dqdPE3);
bproc.minv_block_in_R6_C3_dqdPE3(minv_block_in_R6_C3_dqdPE3);
bproc.minv_block_in_R7_C3_dqdPE3(minv_block_in_R7_C3_dqdPE3);

bproc.minv_block_in_R1_C4_dqdPE3(minv_block_in_R1_C4_dqdPE3);
bproc.minv_block_in_R2_C4_dqdPE3(minv_block_in_R2_C4_dqdPE3);
bproc.minv_block_in_R3_C4_dqdPE3(minv_block_in_R3_C4_dqdPE3);
bproc.minv_block_in_R4_C4_dqdPE3(minv_block_in_R4_C4_dqdPE3);
bproc.minv_block_in_R5_C4_dqdPE3(minv_block_in_R5_C4_dqdPE3);
bproc.minv_block_in_R6_C4_dqdPE3(minv_block_in_R6_C4_dqdPE3);
bproc.minv_block_in_R7_C4_dqdPE3(minv_block_in_R7_C4_dqdPE3);

bproc.minv_block_in_R1_C5_dqdPE3(minv_block_in_R1_C5_dqdPE3);
bproc.minv_block_in_R2_C5_dqdPE3(minv_block_in_R2_C5_dqdPE3);
bproc.minv_block_in_R3_C5_dqdPE3(minv_block_in_R3_C5_dqdPE3);
bproc.minv_block_in_R4_C5_dqdPE3(minv_block_in_R4_C5_dqdPE3);
bproc.minv_block_in_R5_C5_dqdPE3(minv_block_in_R5_C5_dqdPE3);
bproc.minv_block_in_R6_C5_dqdPE3(minv_block_in_R6_C5_dqdPE3);
bproc.minv_block_in_R7_C5_dqdPE3(minv_block_in_R7_C5_dqdPE3);

bproc.minv_block_in_R1_C6_dqdPE3(minv_block_in_R1_C6_dqdPE3);
bproc.minv_block_in_R2_C6_dqdPE3(minv_block_in_R2_C6_dqdPE3);
bproc.minv_block_in_R3_C6_dqdPE3(minv_block_in_R3_C6_dqdPE3);
bproc.minv_block_in_R4_C6_dqdPE3(minv_block_in_R4_C6_dqdPE3);
bproc.minv_block_in_R5_C6_dqdPE3(minv_block_in_R5_C6_dqdPE3);
bproc.minv_block_in_R6_C6_dqdPE3(minv_block_in_R6_C6_dqdPE3);
bproc.minv_block_in_R7_C6_dqdPE3(minv_block_in_R7_C6_dqdPE3);

bproc.minv_block_in_R1_C7_dqdPE3(minv_block_in_R1_C7_dqdPE3);
bproc.minv_block_in_R2_C7_dqdPE3(minv_block_in_R2_C7_dqdPE3);
bproc.minv_block_in_R3_C7_dqdPE3(minv_block_in_R3_C7_dqdPE3);
bproc.minv_block_in_R4_C7_dqdPE3(minv_block_in_R4_C7_dqdPE3);
bproc.minv_block_in_R5_C7_dqdPE3(minv_block_in_R5_C7_dqdPE3);
bproc.minv_block_in_R6_C7_dqdPE3(minv_block_in_R6_C7_dqdPE3);
bproc.minv_block_in_R7_C7_dqdPE3(minv_block_in_R7_C7_dqdPE3);

bproc.dtau_vec_in_R1_dqdPE3(dtau_vec_in_R1_dqdPE3);
bproc.dtau_vec_in_R2_dqdPE3(dtau_vec_in_R2_dqdPE3);
bproc.dtau_vec_in_R3_dqdPE3(dtau_vec_in_R3_dqdPE3);
bproc.dtau_vec_in_R4_dqdPE3(dtau_vec_in_R4_dqdPE3);
bproc.dtau_vec_in_R5_dqdPE3(dtau_vec_in_R5_dqdPE3);
bproc.dtau_vec_in_R6_dqdPE3(dtau_vec_in_R6_dqdPE3);
bproc.dtau_vec_in_R7_dqdPE3(dtau_vec_in_R7_dqdPE3);

bproc.minv_block_in_R1_C1_dqdPE4(minv_block_in_R1_C1_dqdPE4);
bproc.minv_block_in_R2_C1_dqdPE4(minv_block_in_R2_C1_dqdPE4);
bproc.minv_block_in_R3_C1_dqdPE4(minv_block_in_R3_C1_dqdPE4);
bproc.minv_block_in_R4_C1_dqdPE4(minv_block_in_R4_C1_dqdPE4);
bproc.minv_block_in_R5_C1_dqdPE4(minv_block_in_R5_C1_dqdPE4);
bproc.minv_block_in_R6_C1_dqdPE4(minv_block_in_R6_C1_dqdPE4);
bproc.minv_block_in_R7_C1_dqdPE4(minv_block_in_R7_C1_dqdPE4);

bproc.minv_block_in_R1_C2_dqdPE4(minv_block_in_R1_C2_dqdPE4);
bproc.minv_block_in_R2_C2_dqdPE4(minv_block_in_R2_C2_dqdPE4);
bproc.minv_block_in_R3_C2_dqdPE4(minv_block_in_R3_C2_dqdPE4);
bproc.minv_block_in_R4_C2_dqdPE4(minv_block_in_R4_C2_dqdPE4);
bproc.minv_block_in_R5_C2_dqdPE4(minv_block_in_R5_C2_dqdPE4);
bproc.minv_block_in_R6_C2_dqdPE4(minv_block_in_R6_C2_dqdPE4);
bproc.minv_block_in_R7_C2_dqdPE4(minv_block_in_R7_C2_dqdPE4);

bproc.minv_block_in_R1_C3_dqdPE4(minv_block_in_R1_C3_dqdPE4);
bproc.minv_block_in_R2_C3_dqdPE4(minv_block_in_R2_C3_dqdPE4);
bproc.minv_block_in_R3_C3_dqdPE4(minv_block_in_R3_C3_dqdPE4);
bproc.minv_block_in_R4_C3_dqdPE4(minv_block_in_R4_C3_dqdPE4);
bproc.minv_block_in_R5_C3_dqdPE4(minv_block_in_R5_C3_dqdPE4);
bproc.minv_block_in_R6_C3_dqdPE4(minv_block_in_R6_C3_dqdPE4);
bproc.minv_block_in_R7_C3_dqdPE4(minv_block_in_R7_C3_dqdPE4);

bproc.minv_block_in_R1_C4_dqdPE4(minv_block_in_R1_C4_dqdPE4);
bproc.minv_block_in_R2_C4_dqdPE4(minv_block_in_R2_C4_dqdPE4);
bproc.minv_block_in_R3_C4_dqdPE4(minv_block_in_R3_C4_dqdPE4);
bproc.minv_block_in_R4_C4_dqdPE4(minv_block_in_R4_C4_dqdPE4);
bproc.minv_block_in_R5_C4_dqdPE4(minv_block_in_R5_C4_dqdPE4);
bproc.minv_block_in_R6_C4_dqdPE4(minv_block_in_R6_C4_dqdPE4);
bproc.minv_block_in_R7_C4_dqdPE4(minv_block_in_R7_C4_dqdPE4);

bproc.minv_block_in_R1_C5_dqdPE4(minv_block_in_R1_C5_dqdPE4);
bproc.minv_block_in_R2_C5_dqdPE4(minv_block_in_R2_C5_dqdPE4);
bproc.minv_block_in_R3_C5_dqdPE4(minv_block_in_R3_C5_dqdPE4);
bproc.minv_block_in_R4_C5_dqdPE4(minv_block_in_R4_C5_dqdPE4);
bproc.minv_block_in_R5_C5_dqdPE4(minv_block_in_R5_C5_dqdPE4);
bproc.minv_block_in_R6_C5_dqdPE4(minv_block_in_R6_C5_dqdPE4);
bproc.minv_block_in_R7_C5_dqdPE4(minv_block_in_R7_C5_dqdPE4);

bproc.minv_block_in_R1_C6_dqdPE4(minv_block_in_R1_C6_dqdPE4);
bproc.minv_block_in_R2_C6_dqdPE4(minv_block_in_R2_C6_dqdPE4);
bproc.minv_block_in_R3_C6_dqdPE4(minv_block_in_R3_C6_dqdPE4);
bproc.minv_block_in_R4_C6_dqdPE4(minv_block_in_R4_C6_dqdPE4);
bproc.minv_block_in_R5_C6_dqdPE4(minv_block_in_R5_C6_dqdPE4);
bproc.minv_block_in_R6_C6_dqdPE4(minv_block_in_R6_C6_dqdPE4);
bproc.minv_block_in_R7_C6_dqdPE4(minv_block_in_R7_C6_dqdPE4);

bproc.minv_block_in_R1_C7_dqdPE4(minv_block_in_R1_C7_dqdPE4);
bproc.minv_block_in_R2_C7_dqdPE4(minv_block_in_R2_C7_dqdPE4);
bproc.minv_block_in_R3_C7_dqdPE4(minv_block_in_R3_C7_dqdPE4);
bproc.minv_block_in_R4_C7_dqdPE4(minv_block_in_R4_C7_dqdPE4);
bproc.minv_block_in_R5_C7_dqdPE4(minv_block_in_R5_C7_dqdPE4);
bproc.minv_block_in_R6_C7_dqdPE4(minv_block_in_R6_C7_dqdPE4);
bproc.minv_block_in_R7_C7_dqdPE4(minv_block_in_R7_C7_dqdPE4);

bproc.dtau_vec_in_R1_dqdPE4(dtau_vec_in_R1_dqdPE4);
bproc.dtau_vec_in_R2_dqdPE4(dtau_vec_in_R2_dqdPE4);
bproc.dtau_vec_in_R3_dqdPE4(dtau_vec_in_R3_dqdPE4);
bproc.dtau_vec_in_R4_dqdPE4(dtau_vec_in_R4_dqdPE4);
bproc.dtau_vec_in_R5_dqdPE4(dtau_vec_in_R5_dqdPE4);
bproc.dtau_vec_in_R6_dqdPE4(dtau_vec_in_R6_dqdPE4);
bproc.dtau_vec_in_R7_dqdPE4(dtau_vec_in_R7_dqdPE4);

bproc.minv_block_in_R1_C1_dqdPE5(minv_block_in_R1_C1_dqdPE5);
bproc.minv_block_in_R2_C1_dqdPE5(minv_block_in_R2_C1_dqdPE5);
bproc.minv_block_in_R3_C1_dqdPE5(minv_block_in_R3_C1_dqdPE5);
bproc.minv_block_in_R4_C1_dqdPE5(minv_block_in_R4_C1_dqdPE5);
bproc.minv_block_in_R5_C1_dqdPE5(minv_block_in_R5_C1_dqdPE5);
bproc.minv_block_in_R6_C1_dqdPE5(minv_block_in_R6_C1_dqdPE5);
bproc.minv_block_in_R7_C1_dqdPE5(minv_block_in_R7_C1_dqdPE5);

bproc.minv_block_in_R1_C2_dqdPE5(minv_block_in_R1_C2_dqdPE5);
bproc.minv_block_in_R2_C2_dqdPE5(minv_block_in_R2_C2_dqdPE5);
bproc.minv_block_in_R3_C2_dqdPE5(minv_block_in_R3_C2_dqdPE5);
bproc.minv_block_in_R4_C2_dqdPE5(minv_block_in_R4_C2_dqdPE5);
bproc.minv_block_in_R5_C2_dqdPE5(minv_block_in_R5_C2_dqdPE5);
bproc.minv_block_in_R6_C2_dqdPE5(minv_block_in_R6_C2_dqdPE5);
bproc.minv_block_in_R7_C2_dqdPE5(minv_block_in_R7_C2_dqdPE5);

bproc.minv_block_in_R1_C3_dqdPE5(minv_block_in_R1_C3_dqdPE5);
bproc.minv_block_in_R2_C3_dqdPE5(minv_block_in_R2_C3_dqdPE5);
bproc.minv_block_in_R3_C3_dqdPE5(minv_block_in_R3_C3_dqdPE5);
bproc.minv_block_in_R4_C3_dqdPE5(minv_block_in_R4_C3_dqdPE5);
bproc.minv_block_in_R5_C3_dqdPE5(minv_block_in_R5_C3_dqdPE5);
bproc.minv_block_in_R6_C3_dqdPE5(minv_block_in_R6_C3_dqdPE5);
bproc.minv_block_in_R7_C3_dqdPE5(minv_block_in_R7_C3_dqdPE5);

bproc.minv_block_in_R1_C4_dqdPE5(minv_block_in_R1_C4_dqdPE5);
bproc.minv_block_in_R2_C4_dqdPE5(minv_block_in_R2_C4_dqdPE5);
bproc.minv_block_in_R3_C4_dqdPE5(minv_block_in_R3_C4_dqdPE5);
bproc.minv_block_in_R4_C4_dqdPE5(minv_block_in_R4_C4_dqdPE5);
bproc.minv_block_in_R5_C4_dqdPE5(minv_block_in_R5_C4_dqdPE5);
bproc.minv_block_in_R6_C4_dqdPE5(minv_block_in_R6_C4_dqdPE5);
bproc.minv_block_in_R7_C4_dqdPE5(minv_block_in_R7_C4_dqdPE5);

bproc.minv_block_in_R1_C5_dqdPE5(minv_block_in_R1_C5_dqdPE5);
bproc.minv_block_in_R2_C5_dqdPE5(minv_block_in_R2_C5_dqdPE5);
bproc.minv_block_in_R3_C5_dqdPE5(minv_block_in_R3_C5_dqdPE5);
bproc.minv_block_in_R4_C5_dqdPE5(minv_block_in_R4_C5_dqdPE5);
bproc.minv_block_in_R5_C5_dqdPE5(minv_block_in_R5_C5_dqdPE5);
bproc.minv_block_in_R6_C5_dqdPE5(minv_block_in_R6_C5_dqdPE5);
bproc.minv_block_in_R7_C5_dqdPE5(minv_block_in_R7_C5_dqdPE5);

bproc.minv_block_in_R1_C6_dqdPE5(minv_block_in_R1_C6_dqdPE5);
bproc.minv_block_in_R2_C6_dqdPE5(minv_block_in_R2_C6_dqdPE5);
bproc.minv_block_in_R3_C6_dqdPE5(minv_block_in_R3_C6_dqdPE5);
bproc.minv_block_in_R4_C6_dqdPE5(minv_block_in_R4_C6_dqdPE5);
bproc.minv_block_in_R5_C6_dqdPE5(minv_block_in_R5_C6_dqdPE5);
bproc.minv_block_in_R6_C6_dqdPE5(minv_block_in_R6_C6_dqdPE5);
bproc.minv_block_in_R7_C6_dqdPE5(minv_block_in_R7_C6_dqdPE5);

bproc.minv_block_in_R1_C7_dqdPE5(minv_block_in_R1_C7_dqdPE5);
bproc.minv_block_in_R2_C7_dqdPE5(minv_block_in_R2_C7_dqdPE5);
bproc.minv_block_in_R3_C7_dqdPE5(minv_block_in_R3_C7_dqdPE5);
bproc.minv_block_in_R4_C7_dqdPE5(minv_block_in_R4_C7_dqdPE5);
bproc.minv_block_in_R5_C7_dqdPE5(minv_block_in_R5_C7_dqdPE5);
bproc.minv_block_in_R6_C7_dqdPE5(minv_block_in_R6_C7_dqdPE5);
bproc.minv_block_in_R7_C7_dqdPE5(minv_block_in_R7_C7_dqdPE5);

bproc.dtau_vec_in_R1_dqdPE5(dtau_vec_in_R1_dqdPE5);
bproc.dtau_vec_in_R2_dqdPE5(dtau_vec_in_R2_dqdPE5);
bproc.dtau_vec_in_R3_dqdPE5(dtau_vec_in_R3_dqdPE5);
bproc.dtau_vec_in_R4_dqdPE5(dtau_vec_in_R4_dqdPE5);
bproc.dtau_vec_in_R5_dqdPE5(dtau_vec_in_R5_dqdPE5);
bproc.dtau_vec_in_R6_dqdPE5(dtau_vec_in_R6_dqdPE5);
bproc.dtau_vec_in_R7_dqdPE5(dtau_vec_in_R7_dqdPE5);

bproc.minv_block_in_R1_C1_dqdPE6(minv_block_in_R1_C1_dqdPE6);
bproc.minv_block_in_R2_C1_dqdPE6(minv_block_in_R2_C1_dqdPE6);
bproc.minv_block_in_R3_C1_dqdPE6(minv_block_in_R3_C1_dqdPE6);
bproc.minv_block_in_R4_C1_dqdPE6(minv_block_in_R4_C1_dqdPE6);
bproc.minv_block_in_R5_C1_dqdPE6(minv_block_in_R5_C1_dqdPE6);
bproc.minv_block_in_R6_C1_dqdPE6(minv_block_in_R6_C1_dqdPE6);
bproc.minv_block_in_R7_C1_dqdPE6(minv_block_in_R7_C1_dqdPE6);

bproc.minv_block_in_R1_C2_dqdPE6(minv_block_in_R1_C2_dqdPE6);
bproc.minv_block_in_R2_C2_dqdPE6(minv_block_in_R2_C2_dqdPE6);
bproc.minv_block_in_R3_C2_dqdPE6(minv_block_in_R3_C2_dqdPE6);
bproc.minv_block_in_R4_C2_dqdPE6(minv_block_in_R4_C2_dqdPE6);
bproc.minv_block_in_R5_C2_dqdPE6(minv_block_in_R5_C2_dqdPE6);
bproc.minv_block_in_R6_C2_dqdPE6(minv_block_in_R6_C2_dqdPE6);
bproc.minv_block_in_R7_C2_dqdPE6(minv_block_in_R7_C2_dqdPE6);

bproc.minv_block_in_R1_C3_dqdPE6(minv_block_in_R1_C3_dqdPE6);
bproc.minv_block_in_R2_C3_dqdPE6(minv_block_in_R2_C3_dqdPE6);
bproc.minv_block_in_R3_C3_dqdPE6(minv_block_in_R3_C3_dqdPE6);
bproc.minv_block_in_R4_C3_dqdPE6(minv_block_in_R4_C3_dqdPE6);
bproc.minv_block_in_R5_C3_dqdPE6(minv_block_in_R5_C3_dqdPE6);
bproc.minv_block_in_R6_C3_dqdPE6(minv_block_in_R6_C3_dqdPE6);
bproc.minv_block_in_R7_C3_dqdPE6(minv_block_in_R7_C3_dqdPE6);

bproc.minv_block_in_R1_C4_dqdPE6(minv_block_in_R1_C4_dqdPE6);
bproc.minv_block_in_R2_C4_dqdPE6(minv_block_in_R2_C4_dqdPE6);
bproc.minv_block_in_R3_C4_dqdPE6(minv_block_in_R3_C4_dqdPE6);
bproc.minv_block_in_R4_C4_dqdPE6(minv_block_in_R4_C4_dqdPE6);
bproc.minv_block_in_R5_C4_dqdPE6(minv_block_in_R5_C4_dqdPE6);
bproc.minv_block_in_R6_C4_dqdPE6(minv_block_in_R6_C4_dqdPE6);
bproc.minv_block_in_R7_C4_dqdPE6(minv_block_in_R7_C4_dqdPE6);

bproc.minv_block_in_R1_C5_dqdPE6(minv_block_in_R1_C5_dqdPE6);
bproc.minv_block_in_R2_C5_dqdPE6(minv_block_in_R2_C5_dqdPE6);
bproc.minv_block_in_R3_C5_dqdPE6(minv_block_in_R3_C5_dqdPE6);
bproc.minv_block_in_R4_C5_dqdPE6(minv_block_in_R4_C5_dqdPE6);
bproc.minv_block_in_R5_C5_dqdPE6(minv_block_in_R5_C5_dqdPE6);
bproc.minv_block_in_R6_C5_dqdPE6(minv_block_in_R6_C5_dqdPE6);
bproc.minv_block_in_R7_C5_dqdPE6(minv_block_in_R7_C5_dqdPE6);

bproc.minv_block_in_R1_C6_dqdPE6(minv_block_in_R1_C6_dqdPE6);
bproc.minv_block_in_R2_C6_dqdPE6(minv_block_in_R2_C6_dqdPE6);
bproc.minv_block_in_R3_C6_dqdPE6(minv_block_in_R3_C6_dqdPE6);
bproc.minv_block_in_R4_C6_dqdPE6(minv_block_in_R4_C6_dqdPE6);
bproc.minv_block_in_R5_C6_dqdPE6(minv_block_in_R5_C6_dqdPE6);
bproc.minv_block_in_R6_C6_dqdPE6(minv_block_in_R6_C6_dqdPE6);
bproc.minv_block_in_R7_C6_dqdPE6(minv_block_in_R7_C6_dqdPE6);

bproc.minv_block_in_R1_C7_dqdPE6(minv_block_in_R1_C7_dqdPE6);
bproc.minv_block_in_R2_C7_dqdPE6(minv_block_in_R2_C7_dqdPE6);
bproc.minv_block_in_R3_C7_dqdPE6(minv_block_in_R3_C7_dqdPE6);
bproc.minv_block_in_R4_C7_dqdPE6(minv_block_in_R4_C7_dqdPE6);
bproc.minv_block_in_R5_C7_dqdPE6(minv_block_in_R5_C7_dqdPE6);
bproc.minv_block_in_R6_C7_dqdPE6(minv_block_in_R6_C7_dqdPE6);
bproc.minv_block_in_R7_C7_dqdPE6(minv_block_in_R7_C7_dqdPE6);

bproc.dtau_vec_in_R1_dqdPE6(dtau_vec_in_R1_dqdPE6);
bproc.dtau_vec_in_R2_dqdPE6(dtau_vec_in_R2_dqdPE6);
bproc.dtau_vec_in_R3_dqdPE6(dtau_vec_in_R3_dqdPE6);
bproc.dtau_vec_in_R4_dqdPE6(dtau_vec_in_R4_dqdPE6);
bproc.dtau_vec_in_R5_dqdPE6(dtau_vec_in_R5_dqdPE6);
bproc.dtau_vec_in_R6_dqdPE6(dtau_vec_in_R6_dqdPE6);
bproc.dtau_vec_in_R7_dqdPE6(dtau_vec_in_R7_dqdPE6);

bproc.minv_block_in_R1_C1_dqdPE7(minv_block_in_R1_C1_dqdPE7);
bproc.minv_block_in_R2_C1_dqdPE7(minv_block_in_R2_C1_dqdPE7);
bproc.minv_block_in_R3_C1_dqdPE7(minv_block_in_R3_C1_dqdPE7);
bproc.minv_block_in_R4_C1_dqdPE7(minv_block_in_R4_C1_dqdPE7);
bproc.minv_block_in_R5_C1_dqdPE7(minv_block_in_R5_C1_dqdPE7);
bproc.minv_block_in_R6_C1_dqdPE7(minv_block_in_R6_C1_dqdPE7);
bproc.minv_block_in_R7_C1_dqdPE7(minv_block_in_R7_C1_dqdPE7);

bproc.minv_block_in_R1_C2_dqdPE7(minv_block_in_R1_C2_dqdPE7);
bproc.minv_block_in_R2_C2_dqdPE7(minv_block_in_R2_C2_dqdPE7);
bproc.minv_block_in_R3_C2_dqdPE7(minv_block_in_R3_C2_dqdPE7);
bproc.minv_block_in_R4_C2_dqdPE7(minv_block_in_R4_C2_dqdPE7);
bproc.minv_block_in_R5_C2_dqdPE7(minv_block_in_R5_C2_dqdPE7);
bproc.minv_block_in_R6_C2_dqdPE7(minv_block_in_R6_C2_dqdPE7);
bproc.minv_block_in_R7_C2_dqdPE7(minv_block_in_R7_C2_dqdPE7);

bproc.minv_block_in_R1_C3_dqdPE7(minv_block_in_R1_C3_dqdPE7);
bproc.minv_block_in_R2_C3_dqdPE7(minv_block_in_R2_C3_dqdPE7);
bproc.minv_block_in_R3_C3_dqdPE7(minv_block_in_R3_C3_dqdPE7);
bproc.minv_block_in_R4_C3_dqdPE7(minv_block_in_R4_C3_dqdPE7);
bproc.minv_block_in_R5_C3_dqdPE7(minv_block_in_R5_C3_dqdPE7);
bproc.minv_block_in_R6_C3_dqdPE7(minv_block_in_R6_C3_dqdPE7);
bproc.minv_block_in_R7_C3_dqdPE7(minv_block_in_R7_C3_dqdPE7);

bproc.minv_block_in_R1_C4_dqdPE7(minv_block_in_R1_C4_dqdPE7);
bproc.minv_block_in_R2_C4_dqdPE7(minv_block_in_R2_C4_dqdPE7);
bproc.minv_block_in_R3_C4_dqdPE7(minv_block_in_R3_C4_dqdPE7);
bproc.minv_block_in_R4_C4_dqdPE7(minv_block_in_R4_C4_dqdPE7);
bproc.minv_block_in_R5_C4_dqdPE7(minv_block_in_R5_C4_dqdPE7);
bproc.minv_block_in_R6_C4_dqdPE7(minv_block_in_R6_C4_dqdPE7);
bproc.minv_block_in_R7_C4_dqdPE7(minv_block_in_R7_C4_dqdPE7);

bproc.minv_block_in_R1_C5_dqdPE7(minv_block_in_R1_C5_dqdPE7);
bproc.minv_block_in_R2_C5_dqdPE7(minv_block_in_R2_C5_dqdPE7);
bproc.minv_block_in_R3_C5_dqdPE7(minv_block_in_R3_C5_dqdPE7);
bproc.minv_block_in_R4_C5_dqdPE7(minv_block_in_R4_C5_dqdPE7);
bproc.minv_block_in_R5_C5_dqdPE7(minv_block_in_R5_C5_dqdPE7);
bproc.minv_block_in_R6_C5_dqdPE7(minv_block_in_R6_C5_dqdPE7);
bproc.minv_block_in_R7_C5_dqdPE7(minv_block_in_R7_C5_dqdPE7);

bproc.minv_block_in_R1_C6_dqdPE7(minv_block_in_R1_C6_dqdPE7);
bproc.minv_block_in_R2_C6_dqdPE7(minv_block_in_R2_C6_dqdPE7);
bproc.minv_block_in_R3_C6_dqdPE7(minv_block_in_R3_C6_dqdPE7);
bproc.minv_block_in_R4_C6_dqdPE7(minv_block_in_R4_C6_dqdPE7);
bproc.minv_block_in_R5_C6_dqdPE7(minv_block_in_R5_C6_dqdPE7);
bproc.minv_block_in_R6_C6_dqdPE7(minv_block_in_R6_C6_dqdPE7);
bproc.minv_block_in_R7_C6_dqdPE7(minv_block_in_R7_C6_dqdPE7);

bproc.minv_block_in_R1_C7_dqdPE7(minv_block_in_R1_C7_dqdPE7);
bproc.minv_block_in_R2_C7_dqdPE7(minv_block_in_R2_C7_dqdPE7);
bproc.minv_block_in_R3_C7_dqdPE7(minv_block_in_R3_C7_dqdPE7);
bproc.minv_block_in_R4_C7_dqdPE7(minv_block_in_R4_C7_dqdPE7);
bproc.minv_block_in_R5_C7_dqdPE7(minv_block_in_R5_C7_dqdPE7);
bproc.minv_block_in_R6_C7_dqdPE7(minv_block_in_R6_C7_dqdPE7);
bproc.minv_block_in_R7_C7_dqdPE7(minv_block_in_R7_C7_dqdPE7);

bproc.dtau_vec_in_R1_dqdPE7(dtau_vec_in_R1_dqdPE7);
bproc.dtau_vec_in_R2_dqdPE7(dtau_vec_in_R2_dqdPE7);
bproc.dtau_vec_in_R3_dqdPE7(dtau_vec_in_R3_dqdPE7);
bproc.dtau_vec_in_R4_dqdPE7(dtau_vec_in_R4_dqdPE7);
bproc.dtau_vec_in_R5_dqdPE7(dtau_vec_in_R5_dqdPE7);
bproc.dtau_vec_in_R6_dqdPE7(dtau_vec_in_R6_dqdPE7);
bproc.dtau_vec_in_R7_dqdPE7(dtau_vec_in_R7_dqdPE7);

