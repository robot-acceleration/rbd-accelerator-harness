import Clocks::*;
(* always_ready, always_enabled *)
interface BProc;
    (* always_ready *)
    method Action get_data();
    method Action get_data_minv();


    //-------- RNEA INPUTS -----

    method Action link_in_rnea(Bit#(4) v);
    method Action sinq_val_in_rnea(Bit#(32) v);
    method Action cosq_val_in_rnea(Bit#(32) v);

    method Action f_upd_curr_vec_in_AX_rnea(Bit#(32) v);
    method Action f_upd_curr_vec_in_AY_rnea(Bit#(32) v);
    method Action f_upd_curr_vec_in_AZ_rnea(Bit#(32) v);
    method Action f_upd_curr_vec_in_LX_rnea(Bit#(32) v);
    method Action f_upd_curr_vec_in_LY_rnea(Bit#(32) v);
    method Action f_upd_curr_vec_in_LZ_rnea(Bit#(32) v);
    method Action f_prev_vec_in_AX_rnea(Bit#(32) v);
    method Action f_prev_vec_in_AY_rnea(Bit#(32) v);
    method Action f_prev_vec_in_AZ_rnea(Bit#(32) v);
    method Action f_prev_vec_in_LX_rnea(Bit#(32) v);
    method Action f_prev_vec_in_LY_rnea(Bit#(32) v);
    method Action f_prev_vec_in_LZ_rnea(Bit#(32) v);

   //--------------------------

    //-------- DQ AND DQD INPUTS -----

    method Action link_in_dqPE1(Bit#(4) v);
    method Action link_in_dqPE2(Bit#(4) v);
    method Action link_in_dqPE3(Bit#(4) v);
    method Action link_in_dqPE4(Bit#(4) v);
    method Action link_in_dqPE5(Bit#(4) v);
    method Action link_in_dqPE6(Bit#(4) v);
    method Action link_in_dqPE7(Bit#(4) v);
    method Action link_in_dqdPE1(Bit#(4) v);
    method Action link_in_dqdPE2(Bit#(4) v);
    method Action link_in_dqdPE3(Bit#(4) v);
    method Action link_in_dqdPE4(Bit#(4) v);
    method Action link_in_dqdPE5(Bit#(4) v);
    method Action link_in_dqdPE6(Bit#(4) v);
    method Action link_in_dqdPE7(Bit#(4) v);
    method Action derv_in_dqPE1(Bit#(4) v);
    method Action derv_in_dqPE2(Bit#(4) v);
    method Action derv_in_dqPE3(Bit#(4) v);
    method Action derv_in_dqPE4(Bit#(4) v);
    method Action derv_in_dqPE5(Bit#(4) v);
    method Action derv_in_dqPE6(Bit#(4) v);
    method Action derv_in_dqPE7(Bit#(4) v);
    method Action derv_in_dqdPE1(Bit#(4) v);
    method Action derv_in_dqdPE2(Bit#(4) v);
    method Action derv_in_dqdPE3(Bit#(4) v);
    method Action derv_in_dqdPE4(Bit#(4) v);
    method Action derv_in_dqdPE5(Bit#(4) v);
    method Action derv_in_dqdPE6(Bit#(4) v);
    method Action derv_in_dqdPE7(Bit#(4) v);

    method Action sinq_val_in_dqPE1(Bit#(32) v);
    method Action sinq_val_in_dqPE2(Bit#(32) v);
    method Action sinq_val_in_dqPE3(Bit#(32) v);
    method Action sinq_val_in_dqPE4(Bit#(32) v);
    method Action sinq_val_in_dqPE5(Bit#(32) v);
    method Action sinq_val_in_dqPE6(Bit#(32) v);
    method Action sinq_val_in_dqPE7(Bit#(32) v);
    method Action sinq_val_in_dqdPE1(Bit#(32) v);
    method Action sinq_val_in_dqdPE2(Bit#(32) v);
    method Action sinq_val_in_dqdPE3(Bit#(32) v);
    method Action sinq_val_in_dqdPE4(Bit#(32) v);
    method Action sinq_val_in_dqdPE5(Bit#(32) v);
    method Action sinq_val_in_dqdPE6(Bit#(32) v);
    method Action sinq_val_in_dqdPE7(Bit#(32) v);
    method Action cosq_val_in_dqPE1(Bit#(32) v);
    method Action cosq_val_in_dqPE2(Bit#(32) v);
    method Action cosq_val_in_dqPE3(Bit#(32) v);
    method Action cosq_val_in_dqPE4(Bit#(32) v);
    method Action cosq_val_in_dqPE5(Bit#(32) v);
    method Action cosq_val_in_dqPE6(Bit#(32) v);
    method Action cosq_val_in_dqPE7(Bit#(32) v);
    method Action cosq_val_in_dqdPE1(Bit#(32) v);
    method Action cosq_val_in_dqdPE2(Bit#(32) v);
    method Action cosq_val_in_dqdPE3(Bit#(32) v);
    method Action cosq_val_in_dqdPE4(Bit#(32) v);
    method Action cosq_val_in_dqdPE5(Bit#(32) v);
    method Action cosq_val_in_dqdPE6(Bit#(32) v);
    method Action cosq_val_in_dqdPE7(Bit#(32) v);

    method Action f_upd_curr_vec_in_AX_dqPE1(Bit#(32) v);
    method Action f_upd_curr_vec_in_AY_dqPE1(Bit#(32) v);
    method Action f_upd_curr_vec_in_AZ_dqPE1(Bit#(32) v);
    method Action f_upd_curr_vec_in_LX_dqPE1(Bit#(32) v);
    method Action f_upd_curr_vec_in_LY_dqPE1(Bit#(32) v);
    method Action f_upd_curr_vec_in_LZ_dqPE1(Bit#(32) v);
    method Action f_upd_curr_vec_in_AX_dqPE2(Bit#(32) v);
    method Action f_upd_curr_vec_in_AY_dqPE2(Bit#(32) v);
    method Action f_upd_curr_vec_in_AZ_dqPE2(Bit#(32) v);
    method Action f_upd_curr_vec_in_LX_dqPE2(Bit#(32) v);
    method Action f_upd_curr_vec_in_LY_dqPE2(Bit#(32) v);
    method Action f_upd_curr_vec_in_LZ_dqPE2(Bit#(32) v);
    method Action f_upd_curr_vec_in_AX_dqPE3(Bit#(32) v);
    method Action f_upd_curr_vec_in_AY_dqPE3(Bit#(32) v);
    method Action f_upd_curr_vec_in_AZ_dqPE3(Bit#(32) v);
    method Action f_upd_curr_vec_in_LX_dqPE3(Bit#(32) v);
    method Action f_upd_curr_vec_in_LY_dqPE3(Bit#(32) v);
    method Action f_upd_curr_vec_in_LZ_dqPE3(Bit#(32) v);
    method Action f_upd_curr_vec_in_AX_dqPE4(Bit#(32) v);
    method Action f_upd_curr_vec_in_AY_dqPE4(Bit#(32) v);
    method Action f_upd_curr_vec_in_AZ_dqPE4(Bit#(32) v);
    method Action f_upd_curr_vec_in_LX_dqPE4(Bit#(32) v);
    method Action f_upd_curr_vec_in_LY_dqPE4(Bit#(32) v);
    method Action f_upd_curr_vec_in_LZ_dqPE4(Bit#(32) v);
    method Action f_upd_curr_vec_in_AX_dqPE5(Bit#(32) v);
    method Action f_upd_curr_vec_in_AY_dqPE5(Bit#(32) v);
    method Action f_upd_curr_vec_in_AZ_dqPE5(Bit#(32) v);
    method Action f_upd_curr_vec_in_LX_dqPE5(Bit#(32) v);
    method Action f_upd_curr_vec_in_LY_dqPE5(Bit#(32) v);
    method Action f_upd_curr_vec_in_LZ_dqPE5(Bit#(32) v);
    method Action f_upd_curr_vec_in_AX_dqPE6(Bit#(32) v);
    method Action f_upd_curr_vec_in_AY_dqPE6(Bit#(32) v);
    method Action f_upd_curr_vec_in_AZ_dqPE6(Bit#(32) v);
    method Action f_upd_curr_vec_in_LX_dqPE6(Bit#(32) v);
    method Action f_upd_curr_vec_in_LY_dqPE6(Bit#(32) v);
    method Action f_upd_curr_vec_in_LZ_dqPE6(Bit#(32) v);
    method Action f_upd_curr_vec_in_AX_dqPE7(Bit#(32) v);
    method Action f_upd_curr_vec_in_AY_dqPE7(Bit#(32) v);
    method Action f_upd_curr_vec_in_AZ_dqPE7(Bit#(32) v);
    method Action f_upd_curr_vec_in_LX_dqPE7(Bit#(32) v);
    method Action f_upd_curr_vec_in_LY_dqPE7(Bit#(32) v);
    method Action f_upd_curr_vec_in_LZ_dqPE7(Bit#(32) v);
    method Action dfdq_prev_vec_in_AX_dqPE1(Bit#(32) v);
    method Action dfdq_prev_vec_in_AY_dqPE1(Bit#(32) v);
    method Action dfdq_prev_vec_in_AZ_dqPE1(Bit#(32) v);
    method Action dfdq_prev_vec_in_LX_dqPE1(Bit#(32) v);
    method Action dfdq_prev_vec_in_LY_dqPE1(Bit#(32) v);
    method Action dfdq_prev_vec_in_LZ_dqPE1(Bit#(32) v);
    method Action dfdq_prev_vec_in_AX_dqPE2(Bit#(32) v);
    method Action dfdq_prev_vec_in_AY_dqPE2(Bit#(32) v);
    method Action dfdq_prev_vec_in_AZ_dqPE2(Bit#(32) v);
    method Action dfdq_prev_vec_in_LX_dqPE2(Bit#(32) v);
    method Action dfdq_prev_vec_in_LY_dqPE2(Bit#(32) v);
    method Action dfdq_prev_vec_in_LZ_dqPE2(Bit#(32) v);
    method Action dfdq_prev_vec_in_AX_dqPE3(Bit#(32) v);
    method Action dfdq_prev_vec_in_AY_dqPE3(Bit#(32) v);
    method Action dfdq_prev_vec_in_AZ_dqPE3(Bit#(32) v);
    method Action dfdq_prev_vec_in_LX_dqPE3(Bit#(32) v);
    method Action dfdq_prev_vec_in_LY_dqPE3(Bit#(32) v);
    method Action dfdq_prev_vec_in_LZ_dqPE3(Bit#(32) v);
    method Action dfdq_prev_vec_in_AX_dqPE4(Bit#(32) v);
    method Action dfdq_prev_vec_in_AY_dqPE4(Bit#(32) v);
    method Action dfdq_prev_vec_in_AZ_dqPE4(Bit#(32) v);
    method Action dfdq_prev_vec_in_LX_dqPE4(Bit#(32) v);
    method Action dfdq_prev_vec_in_LY_dqPE4(Bit#(32) v);
    method Action dfdq_prev_vec_in_LZ_dqPE4(Bit#(32) v);
    method Action dfdq_prev_vec_in_AX_dqPE5(Bit#(32) v);
    method Action dfdq_prev_vec_in_AY_dqPE5(Bit#(32) v);
    method Action dfdq_prev_vec_in_AZ_dqPE5(Bit#(32) v);
    method Action dfdq_prev_vec_in_LX_dqPE5(Bit#(32) v);
    method Action dfdq_prev_vec_in_LY_dqPE5(Bit#(32) v);
    method Action dfdq_prev_vec_in_LZ_dqPE5(Bit#(32) v);
    method Action dfdq_prev_vec_in_AX_dqPE6(Bit#(32) v);
    method Action dfdq_prev_vec_in_AY_dqPE6(Bit#(32) v);
    method Action dfdq_prev_vec_in_AZ_dqPE6(Bit#(32) v);
    method Action dfdq_prev_vec_in_LX_dqPE6(Bit#(32) v);
    method Action dfdq_prev_vec_in_LY_dqPE6(Bit#(32) v);
    method Action dfdq_prev_vec_in_LZ_dqPE6(Bit#(32) v);
    method Action dfdq_prev_vec_in_AX_dqPE7(Bit#(32) v);
    method Action dfdq_prev_vec_in_AY_dqPE7(Bit#(32) v);
    method Action dfdq_prev_vec_in_AZ_dqPE7(Bit#(32) v);
    method Action dfdq_prev_vec_in_LX_dqPE7(Bit#(32) v);
    method Action dfdq_prev_vec_in_LY_dqPE7(Bit#(32) v);
    method Action dfdq_prev_vec_in_LZ_dqPE7(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AX_dqPE1(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AY_dqPE1(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AZ_dqPE1(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LX_dqPE1(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LY_dqPE1(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LZ_dqPE1(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AX_dqPE2(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AY_dqPE2(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AZ_dqPE2(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LX_dqPE2(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LY_dqPE2(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LZ_dqPE2(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AX_dqPE3(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AY_dqPE3(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AZ_dqPE3(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LX_dqPE3(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LY_dqPE3(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LZ_dqPE3(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AX_dqPE4(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AY_dqPE4(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AZ_dqPE4(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LX_dqPE4(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LY_dqPE4(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LZ_dqPE4(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AX_dqPE5(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AY_dqPE5(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AZ_dqPE5(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LX_dqPE5(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LY_dqPE5(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LZ_dqPE5(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AX_dqPE6(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AY_dqPE6(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AZ_dqPE6(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LX_dqPE6(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LY_dqPE6(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LZ_dqPE6(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AX_dqPE7(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AY_dqPE7(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_AZ_dqPE7(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LX_dqPE7(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LY_dqPE7(Bit#(32) v);
    method Action dfdq_upd_curr_vec_in_LZ_dqPE7(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AX_dqdPE1(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AY_dqdPE1(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AZ_dqdPE1(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LX_dqdPE1(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LY_dqdPE1(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LZ_dqdPE1(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AX_dqdPE2(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AY_dqdPE2(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AZ_dqdPE2(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LX_dqdPE2(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LY_dqdPE2(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LZ_dqdPE2(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AX_dqdPE3(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AY_dqdPE3(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AZ_dqdPE3(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LX_dqdPE3(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LY_dqdPE3(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LZ_dqdPE3(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AX_dqdPE4(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AY_dqdPE4(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AZ_dqdPE4(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LX_dqdPE4(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LY_dqdPE4(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LZ_dqdPE4(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AX_dqdPE5(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AY_dqdPE5(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AZ_dqdPE5(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LX_dqdPE5(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LY_dqdPE5(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LZ_dqdPE5(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AX_dqdPE6(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AY_dqdPE6(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AZ_dqdPE6(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LX_dqdPE6(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LY_dqdPE6(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LZ_dqdPE6(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AX_dqdPE7(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AY_dqdPE7(Bit#(32) v);
    method Action dfdqd_prev_vec_in_AZ_dqdPE7(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LX_dqdPE7(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LY_dqdPE7(Bit#(32) v);
    method Action dfdqd_prev_vec_in_LZ_dqdPE7(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AX_dqdPE1(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AY_dqdPE1(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AZ_dqdPE1(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LX_dqdPE1(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LY_dqdPE1(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LZ_dqdPE1(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AX_dqdPE2(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AY_dqdPE2(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AZ_dqdPE2(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LX_dqdPE2(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LY_dqdPE2(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LZ_dqdPE2(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AX_dqdPE3(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AY_dqdPE3(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AZ_dqdPE3(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LX_dqdPE3(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LY_dqdPE3(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LZ_dqdPE3(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AX_dqdPE4(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AY_dqdPE4(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AZ_dqdPE4(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LX_dqdPE4(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LY_dqdPE4(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LZ_dqdPE4(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AX_dqdPE5(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AY_dqdPE5(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AZ_dqdPE5(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LX_dqdPE5(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LY_dqdPE5(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LZ_dqdPE5(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AX_dqdPE6(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AY_dqdPE6(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AZ_dqdPE6(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LX_dqdPE6(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LY_dqdPE6(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LZ_dqdPE6(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AX_dqdPE7(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AY_dqdPE7(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_AZ_dqdPE7(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LX_dqdPE7(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LY_dqdPE7(Bit#(32) v);
    method Action dfdqd_upd_curr_vec_in_LZ_dqdPE7(Bit#(32) v);

    //-------- MINV EXTERNAL INPUTS -----

    method Action minv_block_in_R1_C1_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R2_C1_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R3_C1_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R4_C1_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R5_C1_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R6_C1_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R7_C1_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R1_C2_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R2_C2_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R3_C2_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R4_C2_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R5_C2_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R6_C2_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R7_C2_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R1_C3_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R2_C3_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R3_C3_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R4_C3_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R5_C3_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R6_C3_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R7_C3_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R1_C4_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R2_C4_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R3_C4_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R4_C4_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R5_C4_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R6_C4_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R7_C4_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R1_C5_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R2_C5_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R3_C5_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R4_C5_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R5_C5_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R6_C5_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R7_C5_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R1_C6_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R2_C6_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R3_C6_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R4_C6_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R5_C6_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R6_C6_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R7_C6_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R1_C7_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R2_C7_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R3_C7_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R4_C7_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R5_C7_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R6_C7_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R7_C7_dqdPE1(Bit#(32) v);
    method Action minv_block_in_R1_C1_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R2_C1_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R3_C1_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R4_C1_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R5_C1_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R6_C1_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R7_C1_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R1_C2_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R2_C2_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R3_C2_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R4_C2_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R5_C2_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R6_C2_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R7_C2_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R1_C3_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R2_C3_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R3_C3_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R4_C3_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R5_C3_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R6_C3_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R7_C3_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R1_C4_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R2_C4_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R3_C4_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R4_C4_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R5_C4_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R6_C4_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R7_C4_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R1_C5_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R2_C5_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R3_C5_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R4_C5_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R5_C5_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R6_C5_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R7_C5_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R1_C6_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R2_C6_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R3_C6_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R4_C6_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R5_C6_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R6_C6_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R7_C6_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R1_C7_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R2_C7_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R3_C7_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R4_C7_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R5_C7_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R6_C7_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R7_C7_dqdPE2(Bit#(32) v);
    method Action minv_block_in_R1_C1_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R2_C1_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R3_C1_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R4_C1_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R5_C1_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R6_C1_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R7_C1_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R1_C2_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R2_C2_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R3_C2_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R4_C2_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R5_C2_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R6_C2_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R7_C2_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R1_C3_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R2_C3_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R3_C3_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R4_C3_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R5_C3_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R6_C3_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R7_C3_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R1_C4_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R2_C4_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R3_C4_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R4_C4_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R5_C4_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R6_C4_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R7_C4_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R1_C5_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R2_C5_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R3_C5_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R4_C5_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R5_C5_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R6_C5_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R7_C5_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R1_C6_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R2_C6_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R3_C6_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R4_C6_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R5_C6_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R6_C6_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R7_C6_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R1_C7_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R2_C7_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R3_C7_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R4_C7_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R5_C7_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R6_C7_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R7_C7_dqdPE3(Bit#(32) v);
    method Action minv_block_in_R1_C1_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R2_C1_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R3_C1_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R4_C1_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R5_C1_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R6_C1_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R7_C1_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R1_C2_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R2_C2_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R3_C2_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R4_C2_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R5_C2_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R6_C2_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R7_C2_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R1_C3_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R2_C3_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R3_C3_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R4_C3_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R5_C3_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R6_C3_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R7_C3_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R1_C4_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R2_C4_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R3_C4_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R4_C4_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R5_C4_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R6_C4_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R7_C4_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R1_C5_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R2_C5_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R3_C5_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R4_C5_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R5_C5_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R6_C5_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R7_C5_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R1_C6_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R2_C6_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R3_C6_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R4_C6_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R5_C6_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R6_C6_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R7_C6_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R1_C7_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R2_C7_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R3_C7_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R4_C7_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R5_C7_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R6_C7_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R7_C7_dqdPE4(Bit#(32) v);
    method Action minv_block_in_R1_C1_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R2_C1_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R3_C1_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R4_C1_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R5_C1_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R6_C1_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R7_C1_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R1_C2_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R2_C2_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R3_C2_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R4_C2_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R5_C2_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R6_C2_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R7_C2_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R1_C3_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R2_C3_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R3_C3_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R4_C3_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R5_C3_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R6_C3_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R7_C3_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R1_C4_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R2_C4_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R3_C4_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R4_C4_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R5_C4_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R6_C4_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R7_C4_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R1_C5_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R2_C5_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R3_C5_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R4_C5_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R5_C5_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R6_C5_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R7_C5_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R1_C6_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R2_C6_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R3_C6_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R4_C6_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R5_C6_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R6_C6_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R7_C6_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R1_C7_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R2_C7_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R3_C7_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R4_C7_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R5_C7_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R6_C7_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R7_C7_dqdPE5(Bit#(32) v);
    method Action minv_block_in_R1_C1_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R2_C1_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R3_C1_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R4_C1_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R5_C1_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R6_C1_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R7_C1_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R1_C2_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R2_C2_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R3_C2_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R4_C2_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R5_C2_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R6_C2_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R7_C2_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R1_C3_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R2_C3_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R3_C3_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R4_C3_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R5_C3_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R6_C3_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R7_C3_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R1_C4_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R2_C4_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R3_C4_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R4_C4_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R5_C4_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R6_C4_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R7_C4_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R1_C5_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R2_C5_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R3_C5_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R4_C5_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R5_C5_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R6_C5_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R7_C5_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R1_C6_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R2_C6_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R3_C6_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R4_C6_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R5_C6_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R6_C6_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R7_C6_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R1_C7_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R2_C7_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R3_C7_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R4_C7_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R5_C7_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R6_C7_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R7_C7_dqdPE6(Bit#(32) v);
    method Action minv_block_in_R1_C1_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R2_C1_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R3_C1_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R4_C1_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R5_C1_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R6_C1_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R7_C1_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R1_C2_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R2_C2_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R3_C2_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R4_C2_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R5_C2_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R6_C2_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R7_C2_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R1_C3_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R2_C3_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R3_C3_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R4_C3_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R5_C3_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R6_C3_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R7_C3_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R1_C4_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R2_C4_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R3_C4_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R4_C4_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R5_C4_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R6_C4_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R7_C4_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R1_C5_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R2_C5_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R3_C5_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R4_C5_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R5_C5_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R6_C5_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R7_C5_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R1_C6_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R2_C6_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R3_C6_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R4_C6_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R5_C6_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R6_C6_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R7_C6_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R1_C7_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R2_C7_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R3_C7_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R4_C7_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R5_C7_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R6_C7_dqdPE7(Bit#(32) v);
    method Action minv_block_in_R7_C7_dqdPE7(Bit#(32) v);
    method Action dtau_vec_in_R1_dqdPE1(Bit#(32) v);
    method Action dtau_vec_in_R2_dqdPE1(Bit#(32) v);
    method Action dtau_vec_in_R3_dqdPE1(Bit#(32) v);
    method Action dtau_vec_in_R4_dqdPE1(Bit#(32) v);
    method Action dtau_vec_in_R5_dqdPE1(Bit#(32) v);
    method Action dtau_vec_in_R6_dqdPE1(Bit#(32) v);
    method Action dtau_vec_in_R7_dqdPE1(Bit#(32) v);
    method Action dtau_vec_in_R1_dqdPE2(Bit#(32) v);
    method Action dtau_vec_in_R2_dqdPE2(Bit#(32) v);
    method Action dtau_vec_in_R3_dqdPE2(Bit#(32) v);
    method Action dtau_vec_in_R4_dqdPE2(Bit#(32) v);
    method Action dtau_vec_in_R5_dqdPE2(Bit#(32) v);
    method Action dtau_vec_in_R6_dqdPE2(Bit#(32) v);
    method Action dtau_vec_in_R7_dqdPE2(Bit#(32) v);
    method Action dtau_vec_in_R1_dqdPE3(Bit#(32) v);
    method Action dtau_vec_in_R2_dqdPE3(Bit#(32) v);
    method Action dtau_vec_in_R3_dqdPE3(Bit#(32) v);
    method Action dtau_vec_in_R4_dqdPE3(Bit#(32) v);
    method Action dtau_vec_in_R5_dqdPE3(Bit#(32) v);
    method Action dtau_vec_in_R6_dqdPE3(Bit#(32) v);
    method Action dtau_vec_in_R7_dqdPE3(Bit#(32) v);
    method Action dtau_vec_in_R1_dqdPE4(Bit#(32) v);
    method Action dtau_vec_in_R2_dqdPE4(Bit#(32) v);
    method Action dtau_vec_in_R3_dqdPE4(Bit#(32) v);
    method Action dtau_vec_in_R4_dqdPE4(Bit#(32) v);
    method Action dtau_vec_in_R5_dqdPE4(Bit#(32) v);
    method Action dtau_vec_in_R6_dqdPE4(Bit#(32) v);
    method Action dtau_vec_in_R7_dqdPE4(Bit#(32) v);
    method Action dtau_vec_in_R1_dqdPE5(Bit#(32) v);
    method Action dtau_vec_in_R2_dqdPE5(Bit#(32) v);
    method Action dtau_vec_in_R3_dqdPE5(Bit#(32) v);
    method Action dtau_vec_in_R4_dqdPE5(Bit#(32) v);
    method Action dtau_vec_in_R5_dqdPE5(Bit#(32) v);
    method Action dtau_vec_in_R6_dqdPE5(Bit#(32) v);
    method Action dtau_vec_in_R7_dqdPE5(Bit#(32) v);
    method Action dtau_vec_in_R1_dqdPE6(Bit#(32) v);
    method Action dtau_vec_in_R2_dqdPE6(Bit#(32) v);
    method Action dtau_vec_in_R3_dqdPE6(Bit#(32) v);
    method Action dtau_vec_in_R4_dqdPE6(Bit#(32) v);
    method Action dtau_vec_in_R5_dqdPE6(Bit#(32) v);
    method Action dtau_vec_in_R6_dqdPE6(Bit#(32) v);
    method Action dtau_vec_in_R7_dqdPE6(Bit#(32) v);
    method Action dtau_vec_in_R1_dqdPE7(Bit#(32) v);
    method Action dtau_vec_in_R2_dqdPE7(Bit#(32) v);
    method Action dtau_vec_in_R3_dqdPE7(Bit#(32) v);
    method Action dtau_vec_in_R4_dqdPE7(Bit#(32) v);
    method Action dtau_vec_in_R5_dqdPE7(Bit#(32) v);
    method Action dtau_vec_in_R6_dqdPE7(Bit#(32) v);
    method Action dtau_vec_in_R7_dqdPE7(Bit#(32) v);

    //--------------------------

    method Bit#(1) output_ready();
    method Bit#(1) output_ready_minv();


    //-------- RNEA OUTPUTS -----

    method Bit#(32) tau_curr_out_rnea();
    method Bit#(32) f_upd_prev_vec_out_AX_rnea();
    method Bit#(32) f_upd_prev_vec_out_AY_rnea();
    method Bit#(32) f_upd_prev_vec_out_AZ_rnea();
    method Bit#(32) f_upd_prev_vec_out_LX_rnea();
    method Bit#(32) f_upd_prev_vec_out_LY_rnea();
    method Bit#(32) f_upd_prev_vec_out_LZ_rnea();

    //-----------------------

    //----------- DQ DQD OUTPUTS -----

    method Bit#(32) dtau_curr_out_dqPE1();
    method Bit#(32) dtau_curr_out_dqPE2();
    method Bit#(32) dtau_curr_out_dqPE3();
    method Bit#(32) dtau_curr_out_dqPE4();
    method Bit#(32) dtau_curr_out_dqPE5();
    method Bit#(32) dtau_curr_out_dqPE6();
    method Bit#(32) dtau_curr_out_dqPE7();
    method Bit#(32) dtau_curr_out_dqdPE1();
    method Bit#(32) dtau_curr_out_dqdPE2();
    method Bit#(32) dtau_curr_out_dqdPE3();
    method Bit#(32) dtau_curr_out_dqdPE4();
    method Bit#(32) dtau_curr_out_dqdPE5();
    method Bit#(32) dtau_curr_out_dqdPE6();
    method Bit#(32) dtau_curr_out_dqdPE7();
    method Bit#(32) dfdq_upd_prev_vec_out_AX_dqPE1();
    method Bit#(32) dfdq_upd_prev_vec_out_AY_dqPE1();
    method Bit#(32) dfdq_upd_prev_vec_out_AZ_dqPE1();
    method Bit#(32) dfdq_upd_prev_vec_out_LX_dqPE1();
    method Bit#(32) dfdq_upd_prev_vec_out_LY_dqPE1();
    method Bit#(32) dfdq_upd_prev_vec_out_LZ_dqPE1();
    method Bit#(32) dfdq_upd_prev_vec_out_AX_dqPE2();
    method Bit#(32) dfdq_upd_prev_vec_out_AY_dqPE2();
    method Bit#(32) dfdq_upd_prev_vec_out_AZ_dqPE2();
    method Bit#(32) dfdq_upd_prev_vec_out_LX_dqPE2();
    method Bit#(32) dfdq_upd_prev_vec_out_LY_dqPE2();
    method Bit#(32) dfdq_upd_prev_vec_out_LZ_dqPE2();
    method Bit#(32) dfdq_upd_prev_vec_out_AX_dqPE3();
    method Bit#(32) dfdq_upd_prev_vec_out_AY_dqPE3();
    method Bit#(32) dfdq_upd_prev_vec_out_AZ_dqPE3();
    method Bit#(32) dfdq_upd_prev_vec_out_LX_dqPE3();
    method Bit#(32) dfdq_upd_prev_vec_out_LY_dqPE3();
    method Bit#(32) dfdq_upd_prev_vec_out_LZ_dqPE3();
    method Bit#(32) dfdq_upd_prev_vec_out_AX_dqPE4();
    method Bit#(32) dfdq_upd_prev_vec_out_AY_dqPE4();
    method Bit#(32) dfdq_upd_prev_vec_out_AZ_dqPE4();
    method Bit#(32) dfdq_upd_prev_vec_out_LX_dqPE4();
    method Bit#(32) dfdq_upd_prev_vec_out_LY_dqPE4();
    method Bit#(32) dfdq_upd_prev_vec_out_LZ_dqPE4();
    method Bit#(32) dfdq_upd_prev_vec_out_AX_dqPE5();
    method Bit#(32) dfdq_upd_prev_vec_out_AY_dqPE5();
    method Bit#(32) dfdq_upd_prev_vec_out_AZ_dqPE5();
    method Bit#(32) dfdq_upd_prev_vec_out_LX_dqPE5();
    method Bit#(32) dfdq_upd_prev_vec_out_LY_dqPE5();
    method Bit#(32) dfdq_upd_prev_vec_out_LZ_dqPE5();
    method Bit#(32) dfdq_upd_prev_vec_out_AX_dqPE6();
    method Bit#(32) dfdq_upd_prev_vec_out_AY_dqPE6();
    method Bit#(32) dfdq_upd_prev_vec_out_AZ_dqPE6();
    method Bit#(32) dfdq_upd_prev_vec_out_LX_dqPE6();
    method Bit#(32) dfdq_upd_prev_vec_out_LY_dqPE6();
    method Bit#(32) dfdq_upd_prev_vec_out_LZ_dqPE6();
    method Bit#(32) dfdq_upd_prev_vec_out_AX_dqPE7();
    method Bit#(32) dfdq_upd_prev_vec_out_AY_dqPE7();
    method Bit#(32) dfdq_upd_prev_vec_out_AZ_dqPE7();
    method Bit#(32) dfdq_upd_prev_vec_out_LX_dqPE7();
    method Bit#(32) dfdq_upd_prev_vec_out_LY_dqPE7();
    method Bit#(32) dfdq_upd_prev_vec_out_LZ_dqPE7();
    method Bit#(32) dfdqd_upd_prev_vec_out_AX_dqdPE1();
    method Bit#(32) dfdqd_upd_prev_vec_out_AY_dqdPE1();
    method Bit#(32) dfdqd_upd_prev_vec_out_AZ_dqdPE1();
    method Bit#(32) dfdqd_upd_prev_vec_out_LX_dqdPE1();
    method Bit#(32) dfdqd_upd_prev_vec_out_LY_dqdPE1();
    method Bit#(32) dfdqd_upd_prev_vec_out_LZ_dqdPE1();
    method Bit#(32) dfdqd_upd_prev_vec_out_AX_dqdPE2();
    method Bit#(32) dfdqd_upd_prev_vec_out_AY_dqdPE2();
    method Bit#(32) dfdqd_upd_prev_vec_out_AZ_dqdPE2();
    method Bit#(32) dfdqd_upd_prev_vec_out_LX_dqdPE2();
    method Bit#(32) dfdqd_upd_prev_vec_out_LY_dqdPE2();
    method Bit#(32) dfdqd_upd_prev_vec_out_LZ_dqdPE2();
    method Bit#(32) dfdqd_upd_prev_vec_out_AX_dqdPE3();
    method Bit#(32) dfdqd_upd_prev_vec_out_AY_dqdPE3();
    method Bit#(32) dfdqd_upd_prev_vec_out_AZ_dqdPE3();
    method Bit#(32) dfdqd_upd_prev_vec_out_LX_dqdPE3();
    method Bit#(32) dfdqd_upd_prev_vec_out_LY_dqdPE3();
    method Bit#(32) dfdqd_upd_prev_vec_out_LZ_dqdPE3();
    method Bit#(32) dfdqd_upd_prev_vec_out_AX_dqdPE4();
    method Bit#(32) dfdqd_upd_prev_vec_out_AY_dqdPE4();
    method Bit#(32) dfdqd_upd_prev_vec_out_AZ_dqdPE4();
    method Bit#(32) dfdqd_upd_prev_vec_out_LX_dqdPE4();
    method Bit#(32) dfdqd_upd_prev_vec_out_LY_dqdPE4();
    method Bit#(32) dfdqd_upd_prev_vec_out_LZ_dqdPE4();
    method Bit#(32) dfdqd_upd_prev_vec_out_AX_dqdPE5();
    method Bit#(32) dfdqd_upd_prev_vec_out_AY_dqdPE5();
    method Bit#(32) dfdqd_upd_prev_vec_out_AZ_dqdPE5();
    method Bit#(32) dfdqd_upd_prev_vec_out_LX_dqdPE5();
    method Bit#(32) dfdqd_upd_prev_vec_out_LY_dqdPE5();
    method Bit#(32) dfdqd_upd_prev_vec_out_LZ_dqdPE5();
    method Bit#(32) dfdqd_upd_prev_vec_out_AX_dqdPE6();
    method Bit#(32) dfdqd_upd_prev_vec_out_AY_dqdPE6();
    method Bit#(32) dfdqd_upd_prev_vec_out_AZ_dqdPE6();
    method Bit#(32) dfdqd_upd_prev_vec_out_LX_dqdPE6();
    method Bit#(32) dfdqd_upd_prev_vec_out_LY_dqdPE6();
    method Bit#(32) dfdqd_upd_prev_vec_out_LZ_dqdPE6();
    method Bit#(32) dfdqd_upd_prev_vec_out_AX_dqdPE7();
    method Bit#(32) dfdqd_upd_prev_vec_out_AY_dqdPE7();
    method Bit#(32) dfdqd_upd_prev_vec_out_AZ_dqdPE7();
    method Bit#(32) dfdqd_upd_prev_vec_out_LX_dqdPE7();
    method Bit#(32) dfdqd_upd_prev_vec_out_LY_dqdPE7();
    method Bit#(32) dfdqd_upd_prev_vec_out_LZ_dqdPE7();

    //----------- MINV EXTERNAL OUTPUTS -----

    method Bit#(32) minv_vec_out_R1_dqdPE1();
    method Bit#(32) minv_vec_out_R2_dqdPE1();
    method Bit#(32) minv_vec_out_R3_dqdPE1();
    method Bit#(32) minv_vec_out_R4_dqdPE1();
    method Bit#(32) minv_vec_out_R5_dqdPE1();
    method Bit#(32) minv_vec_out_R6_dqdPE1();
    method Bit#(32) minv_vec_out_R7_dqdPE1();
    method Bit#(32) minv_vec_out_R1_dqdPE2();
    method Bit#(32) minv_vec_out_R2_dqdPE2();
    method Bit#(32) minv_vec_out_R3_dqdPE2();
    method Bit#(32) minv_vec_out_R4_dqdPE2();
    method Bit#(32) minv_vec_out_R5_dqdPE2();
    method Bit#(32) minv_vec_out_R6_dqdPE2();
    method Bit#(32) minv_vec_out_R7_dqdPE2();
    method Bit#(32) minv_vec_out_R1_dqdPE3();
    method Bit#(32) minv_vec_out_R2_dqdPE3();
    method Bit#(32) minv_vec_out_R3_dqdPE3();
    method Bit#(32) minv_vec_out_R4_dqdPE3();
    method Bit#(32) minv_vec_out_R5_dqdPE3();
    method Bit#(32) minv_vec_out_R6_dqdPE3();
    method Bit#(32) minv_vec_out_R7_dqdPE3();
    method Bit#(32) minv_vec_out_R1_dqdPE4();
    method Bit#(32) minv_vec_out_R2_dqdPE4();
    method Bit#(32) minv_vec_out_R3_dqdPE4();
    method Bit#(32) minv_vec_out_R4_dqdPE4();
    method Bit#(32) minv_vec_out_R5_dqdPE4();
    method Bit#(32) minv_vec_out_R6_dqdPE4();
    method Bit#(32) minv_vec_out_R7_dqdPE4();
    method Bit#(32) minv_vec_out_R1_dqdPE5();
    method Bit#(32) minv_vec_out_R2_dqdPE5();
    method Bit#(32) minv_vec_out_R3_dqdPE5();
    method Bit#(32) minv_vec_out_R4_dqdPE5();
    method Bit#(32) minv_vec_out_R5_dqdPE5();
    method Bit#(32) minv_vec_out_R6_dqdPE5();
    method Bit#(32) minv_vec_out_R7_dqdPE5();
    method Bit#(32) minv_vec_out_R1_dqdPE6();
    method Bit#(32) minv_vec_out_R2_dqdPE6();
    method Bit#(32) minv_vec_out_R3_dqdPE6();
    method Bit#(32) minv_vec_out_R4_dqdPE6();
    method Bit#(32) minv_vec_out_R5_dqdPE6();
    method Bit#(32) minv_vec_out_R6_dqdPE6();
    method Bit#(32) minv_vec_out_R7_dqdPE6();
    method Bit#(32) minv_vec_out_R1_dqdPE7();
    method Bit#(32) minv_vec_out_R2_dqdPE7();
    method Bit#(32) minv_vec_out_R3_dqdPE7();
    method Bit#(32) minv_vec_out_R4_dqdPE7();
    method Bit#(32) minv_vec_out_R5_dqdPE7();
    method Bit#(32) minv_vec_out_R6_dqdPE7();
    method Bit#(32) minv_vec_out_R7_dqdPE7();

endinterface

import "BVI" bproc =
module mkBProc(BProc);
   default_clock clk();
    default_reset rst();
    input_clock (clk) <- exposeCurrentClock; 
    input_reset (reset) <- invertCurrentReset;
    method get_data() enable(get_data);
    method get_data_minv() enable(get_data_minv);


    method link_in_rnea(link_in_rnea) enable((*inhigh*) EN_link_in_rnea) ;
    method sinq_val_in_rnea(sinq_val_in_rnea) enable((*inhigh*) EN_sinq_val_in_rnea) ;
    method cosq_val_in_rnea(cosq_val_in_rnea) enable((*inhigh*) EN_cosq_val_in_rnea) ;

    method f_upd_curr_vec_in_AX_rnea(f_upd_curr_vec_in_AX_rnea) enable((*inhigh*) EN_f_upd_curr_vec_in_AX_rnea) ;
    method f_upd_curr_vec_in_AY_rnea(f_upd_curr_vec_in_AY_rnea) enable((*inhigh*) EN_f_upd_curr_vec_in_AY_rnea) ;
    method f_upd_curr_vec_in_AZ_rnea(f_upd_curr_vec_in_AZ_rnea) enable((*inhigh*) EN_f_upd_curr_vec_in_AZ_rnea) ;
    method f_upd_curr_vec_in_LX_rnea(f_upd_curr_vec_in_LX_rnea) enable((*inhigh*) EN_f_upd_curr_vec_in_LX_rnea) ;
    method f_upd_curr_vec_in_LY_rnea(f_upd_curr_vec_in_LY_rnea) enable((*inhigh*) EN_f_upd_curr_vec_in_LY_rnea) ;
    method f_upd_curr_vec_in_LZ_rnea(f_upd_curr_vec_in_LZ_rnea) enable((*inhigh*) EN_f_upd_curr_vec_in_LZ_rnea) ;
    method f_prev_vec_in_AX_rnea(f_prev_vec_in_AX_rnea) enable((*inhigh*) EN_f_prev_vec_in_AX_rnea) ;
    method f_prev_vec_in_AY_rnea(f_prev_vec_in_AY_rnea) enable((*inhigh*) EN_f_prev_vec_in_AY_rnea) ;
    method f_prev_vec_in_AZ_rnea(f_prev_vec_in_AZ_rnea) enable((*inhigh*) EN_f_prev_vec_in_AZ_rnea) ;
    method f_prev_vec_in_LX_rnea(f_prev_vec_in_LX_rnea) enable((*inhigh*) EN_f_prev_vec_in_LX_rnea) ;
    method f_prev_vec_in_LY_rnea(f_prev_vec_in_LY_rnea) enable((*inhigh*) EN_f_prev_vec_in_LY_rnea) ;
    method f_prev_vec_in_LZ_rnea(f_prev_vec_in_LZ_rnea) enable((*inhigh*) EN_f_prev_vec_in_LZ_rnea) ;

    method link_in_dqPE1(link_in_dqPE1) enable((*inhigh*) EN_link_in_dqPE1) ;
    method link_in_dqPE2(link_in_dqPE2) enable((*inhigh*) EN_link_in_dqPE2) ;
    method link_in_dqPE3(link_in_dqPE3) enable((*inhigh*) EN_link_in_dqPE3) ;
    method link_in_dqPE4(link_in_dqPE4) enable((*inhigh*) EN_link_in_dqPE4) ;
    method link_in_dqPE5(link_in_dqPE5) enable((*inhigh*) EN_link_in_dqPE5) ;
    method link_in_dqPE6(link_in_dqPE6) enable((*inhigh*) EN_link_in_dqPE6) ;
    method link_in_dqPE7(link_in_dqPE7) enable((*inhigh*) EN_link_in_dqPE7) ;
    method link_in_dqdPE1(link_in_dqdPE1) enable((*inhigh*) EN_link_in_dqdPE1) ;
    method link_in_dqdPE2(link_in_dqdPE2) enable((*inhigh*) EN_link_in_dqdPE2) ;
    method link_in_dqdPE3(link_in_dqdPE3) enable((*inhigh*) EN_link_in_dqdPE3) ;
    method link_in_dqdPE4(link_in_dqdPE4) enable((*inhigh*) EN_link_in_dqdPE4) ;
    method link_in_dqdPE5(link_in_dqdPE5) enable((*inhigh*) EN_link_in_dqdPE5) ;
    method link_in_dqdPE6(link_in_dqdPE6) enable((*inhigh*) EN_link_in_dqdPE6) ;
    method link_in_dqdPE7(link_in_dqdPE7) enable((*inhigh*) EN_link_in_dqdPE7) ;
    method derv_in_dqPE1(derv_in_dqPE1) enable((*inhigh*) EN_derv_in_dqPE1) ;
    method derv_in_dqPE2(derv_in_dqPE2) enable((*inhigh*) EN_derv_in_dqPE2) ;
    method derv_in_dqPE3(derv_in_dqPE3) enable((*inhigh*) EN_derv_in_dqPE3) ;
    method derv_in_dqPE4(derv_in_dqPE4) enable((*inhigh*) EN_derv_in_dqPE4) ;
    method derv_in_dqPE5(derv_in_dqPE5) enable((*inhigh*) EN_derv_in_dqPE5) ;
    method derv_in_dqPE6(derv_in_dqPE6) enable((*inhigh*) EN_derv_in_dqPE6) ;
    method derv_in_dqPE7(derv_in_dqPE7) enable((*inhigh*) EN_derv_in_dqPE7) ;
    method derv_in_dqdPE1(derv_in_dqdPE1) enable((*inhigh*) EN_derv_in_dqdPE1) ;
    method derv_in_dqdPE2(derv_in_dqdPE2) enable((*inhigh*) EN_derv_in_dqdPE2) ;
    method derv_in_dqdPE3(derv_in_dqdPE3) enable((*inhigh*) EN_derv_in_dqdPE3) ;
    method derv_in_dqdPE4(derv_in_dqdPE4) enable((*inhigh*) EN_derv_in_dqdPE4) ;
    method derv_in_dqdPE5(derv_in_dqdPE5) enable((*inhigh*) EN_derv_in_dqdPE5) ;
    method derv_in_dqdPE6(derv_in_dqdPE6) enable((*inhigh*) EN_derv_in_dqdPE6) ;
    method derv_in_dqdPE7(derv_in_dqdPE7) enable((*inhigh*) EN_derv_in_dqdPE7) ;

    method sinq_val_in_dqPE1(sinq_val_in_dqPE1) enable((*inhigh*) EN_sinq_val_in_dqPE1) ;
    method sinq_val_in_dqPE2(sinq_val_in_dqPE2) enable((*inhigh*) EN_sinq_val_in_dqPE2) ;
    method sinq_val_in_dqPE3(sinq_val_in_dqPE3) enable((*inhigh*) EN_sinq_val_in_dqPE3) ;
    method sinq_val_in_dqPE4(sinq_val_in_dqPE4) enable((*inhigh*) EN_sinq_val_in_dqPE4) ;
    method sinq_val_in_dqPE5(sinq_val_in_dqPE5) enable((*inhigh*) EN_sinq_val_in_dqPE5) ;
    method sinq_val_in_dqPE6(sinq_val_in_dqPE6) enable((*inhigh*) EN_sinq_val_in_dqPE6) ;
    method sinq_val_in_dqPE7(sinq_val_in_dqPE7) enable((*inhigh*) EN_sinq_val_in_dqPE7) ;
    method sinq_val_in_dqdPE1(sinq_val_in_dqdPE1) enable((*inhigh*) EN_sinq_val_in_dqdPE1) ;
    method sinq_val_in_dqdPE2(sinq_val_in_dqdPE2) enable((*inhigh*) EN_sinq_val_in_dqdPE2) ;
    method sinq_val_in_dqdPE3(sinq_val_in_dqdPE3) enable((*inhigh*) EN_sinq_val_in_dqdPE3) ;
    method sinq_val_in_dqdPE4(sinq_val_in_dqdPE4) enable((*inhigh*) EN_sinq_val_in_dqdPE4) ;
    method sinq_val_in_dqdPE5(sinq_val_in_dqdPE5) enable((*inhigh*) EN_sinq_val_in_dqdPE5) ;
    method sinq_val_in_dqdPE6(sinq_val_in_dqdPE6) enable((*inhigh*) EN_sinq_val_in_dqdPE6) ;
    method sinq_val_in_dqdPE7(sinq_val_in_dqdPE7) enable((*inhigh*) EN_sinq_val_in_dqdPE7) ;
    method cosq_val_in_dqPE1(cosq_val_in_dqPE1) enable((*inhigh*) EN_cosq_val_in_dqPE1) ;
    method cosq_val_in_dqPE2(cosq_val_in_dqPE2) enable((*inhigh*) EN_cosq_val_in_dqPE2) ;
    method cosq_val_in_dqPE3(cosq_val_in_dqPE3) enable((*inhigh*) EN_cosq_val_in_dqPE3) ;
    method cosq_val_in_dqPE4(cosq_val_in_dqPE4) enable((*inhigh*) EN_cosq_val_in_dqPE4) ;
    method cosq_val_in_dqPE5(cosq_val_in_dqPE5) enable((*inhigh*) EN_cosq_val_in_dqPE5) ;
    method cosq_val_in_dqPE6(cosq_val_in_dqPE6) enable((*inhigh*) EN_cosq_val_in_dqPE6) ;
    method cosq_val_in_dqPE7(cosq_val_in_dqPE7) enable((*inhigh*) EN_cosq_val_in_dqPE7) ;
    method cosq_val_in_dqdPE1(cosq_val_in_dqdPE1) enable((*inhigh*) EN_cosq_val_in_dqdPE1) ;
    method cosq_val_in_dqdPE2(cosq_val_in_dqdPE2) enable((*inhigh*) EN_cosq_val_in_dqdPE2) ;
    method cosq_val_in_dqdPE3(cosq_val_in_dqdPE3) enable((*inhigh*) EN_cosq_val_in_dqdPE3) ;
    method cosq_val_in_dqdPE4(cosq_val_in_dqdPE4) enable((*inhigh*) EN_cosq_val_in_dqdPE4) ;
    method cosq_val_in_dqdPE5(cosq_val_in_dqdPE5) enable((*inhigh*) EN_cosq_val_in_dqdPE5) ;
    method cosq_val_in_dqdPE6(cosq_val_in_dqdPE6) enable((*inhigh*) EN_cosq_val_in_dqdPE6) ;
    method cosq_val_in_dqdPE7(cosq_val_in_dqdPE7) enable((*inhigh*) EN_cosq_val_in_dqdPE7) ;

    method f_upd_curr_vec_in_AX_dqPE1(f_upd_curr_vec_in_AX_dqPE1) enable((*inhigh*) EN_f_upd_curr_vec_in_AX_dqPE1) ;
    method f_upd_curr_vec_in_AY_dqPE1(f_upd_curr_vec_in_AY_dqPE1) enable((*inhigh*) EN_f_upd_curr_vec_in_AY_dqPE1) ;
    method f_upd_curr_vec_in_AZ_dqPE1(f_upd_curr_vec_in_AZ_dqPE1) enable((*inhigh*) EN_f_upd_curr_vec_in_AZ_dqPE1) ;
    method f_upd_curr_vec_in_LX_dqPE1(f_upd_curr_vec_in_LX_dqPE1) enable((*inhigh*) EN_f_upd_curr_vec_in_LX_dqPE1) ;
    method f_upd_curr_vec_in_LY_dqPE1(f_upd_curr_vec_in_LY_dqPE1) enable((*inhigh*) EN_f_upd_curr_vec_in_LY_dqPE1) ;
    method f_upd_curr_vec_in_LZ_dqPE1(f_upd_curr_vec_in_LZ_dqPE1) enable((*inhigh*) EN_f_upd_curr_vec_in_LZ_dqPE1) ;
    method f_upd_curr_vec_in_AX_dqPE2(f_upd_curr_vec_in_AX_dqPE2) enable((*inhigh*) EN_f_upd_curr_vec_in_AX_dqPE2) ;
    method f_upd_curr_vec_in_AY_dqPE2(f_upd_curr_vec_in_AY_dqPE2) enable((*inhigh*) EN_f_upd_curr_vec_in_AY_dqPE2) ;
    method f_upd_curr_vec_in_AZ_dqPE2(f_upd_curr_vec_in_AZ_dqPE2) enable((*inhigh*) EN_f_upd_curr_vec_in_AZ_dqPE2) ;
    method f_upd_curr_vec_in_LX_dqPE2(f_upd_curr_vec_in_LX_dqPE2) enable((*inhigh*) EN_f_upd_curr_vec_in_LX_dqPE2) ;
    method f_upd_curr_vec_in_LY_dqPE2(f_upd_curr_vec_in_LY_dqPE2) enable((*inhigh*) EN_f_upd_curr_vec_in_LY_dqPE2) ;
    method f_upd_curr_vec_in_LZ_dqPE2(f_upd_curr_vec_in_LZ_dqPE2) enable((*inhigh*) EN_f_upd_curr_vec_in_LZ_dqPE2) ;
    method f_upd_curr_vec_in_AX_dqPE3(f_upd_curr_vec_in_AX_dqPE3) enable((*inhigh*) EN_f_upd_curr_vec_in_AX_dqPE3) ;
    method f_upd_curr_vec_in_AY_dqPE3(f_upd_curr_vec_in_AY_dqPE3) enable((*inhigh*) EN_f_upd_curr_vec_in_AY_dqPE3) ;
    method f_upd_curr_vec_in_AZ_dqPE3(f_upd_curr_vec_in_AZ_dqPE3) enable((*inhigh*) EN_f_upd_curr_vec_in_AZ_dqPE3) ;
    method f_upd_curr_vec_in_LX_dqPE3(f_upd_curr_vec_in_LX_dqPE3) enable((*inhigh*) EN_f_upd_curr_vec_in_LX_dqPE3) ;
    method f_upd_curr_vec_in_LY_dqPE3(f_upd_curr_vec_in_LY_dqPE3) enable((*inhigh*) EN_f_upd_curr_vec_in_LY_dqPE3) ;
    method f_upd_curr_vec_in_LZ_dqPE3(f_upd_curr_vec_in_LZ_dqPE3) enable((*inhigh*) EN_f_upd_curr_vec_in_LZ_dqPE3) ;
    method f_upd_curr_vec_in_AX_dqPE4(f_upd_curr_vec_in_AX_dqPE4) enable((*inhigh*) EN_f_upd_curr_vec_in_AX_dqPE4) ;
    method f_upd_curr_vec_in_AY_dqPE4(f_upd_curr_vec_in_AY_dqPE4) enable((*inhigh*) EN_f_upd_curr_vec_in_AY_dqPE4) ;
    method f_upd_curr_vec_in_AZ_dqPE4(f_upd_curr_vec_in_AZ_dqPE4) enable((*inhigh*) EN_f_upd_curr_vec_in_AZ_dqPE4) ;
    method f_upd_curr_vec_in_LX_dqPE4(f_upd_curr_vec_in_LX_dqPE4) enable((*inhigh*) EN_f_upd_curr_vec_in_LX_dqPE4) ;
    method f_upd_curr_vec_in_LY_dqPE4(f_upd_curr_vec_in_LY_dqPE4) enable((*inhigh*) EN_f_upd_curr_vec_in_LY_dqPE4) ;
    method f_upd_curr_vec_in_LZ_dqPE4(f_upd_curr_vec_in_LZ_dqPE4) enable((*inhigh*) EN_f_upd_curr_vec_in_LZ_dqPE4) ;
    method f_upd_curr_vec_in_AX_dqPE5(f_upd_curr_vec_in_AX_dqPE5) enable((*inhigh*) EN_f_upd_curr_vec_in_AX_dqPE5) ;
    method f_upd_curr_vec_in_AY_dqPE5(f_upd_curr_vec_in_AY_dqPE5) enable((*inhigh*) EN_f_upd_curr_vec_in_AY_dqPE5) ;
    method f_upd_curr_vec_in_AZ_dqPE5(f_upd_curr_vec_in_AZ_dqPE5) enable((*inhigh*) EN_f_upd_curr_vec_in_AZ_dqPE5) ;
    method f_upd_curr_vec_in_LX_dqPE5(f_upd_curr_vec_in_LX_dqPE5) enable((*inhigh*) EN_f_upd_curr_vec_in_LX_dqPE5) ;
    method f_upd_curr_vec_in_LY_dqPE5(f_upd_curr_vec_in_LY_dqPE5) enable((*inhigh*) EN_f_upd_curr_vec_in_LY_dqPE5) ;
    method f_upd_curr_vec_in_LZ_dqPE5(f_upd_curr_vec_in_LZ_dqPE5) enable((*inhigh*) EN_f_upd_curr_vec_in_LZ_dqPE5) ;
    method f_upd_curr_vec_in_AX_dqPE6(f_upd_curr_vec_in_AX_dqPE6) enable((*inhigh*) EN_f_upd_curr_vec_in_AX_dqPE6) ;
    method f_upd_curr_vec_in_AY_dqPE6(f_upd_curr_vec_in_AY_dqPE6) enable((*inhigh*) EN_f_upd_curr_vec_in_AY_dqPE6) ;
    method f_upd_curr_vec_in_AZ_dqPE6(f_upd_curr_vec_in_AZ_dqPE6) enable((*inhigh*) EN_f_upd_curr_vec_in_AZ_dqPE6) ;
    method f_upd_curr_vec_in_LX_dqPE6(f_upd_curr_vec_in_LX_dqPE6) enable((*inhigh*) EN_f_upd_curr_vec_in_LX_dqPE6) ;
    method f_upd_curr_vec_in_LY_dqPE6(f_upd_curr_vec_in_LY_dqPE6) enable((*inhigh*) EN_f_upd_curr_vec_in_LY_dqPE6) ;
    method f_upd_curr_vec_in_LZ_dqPE6(f_upd_curr_vec_in_LZ_dqPE6) enable((*inhigh*) EN_f_upd_curr_vec_in_LZ_dqPE6) ;
    method f_upd_curr_vec_in_AX_dqPE7(f_upd_curr_vec_in_AX_dqPE7) enable((*inhigh*) EN_f_upd_curr_vec_in_AX_dqPE7) ;
    method f_upd_curr_vec_in_AY_dqPE7(f_upd_curr_vec_in_AY_dqPE7) enable((*inhigh*) EN_f_upd_curr_vec_in_AY_dqPE7) ;
    method f_upd_curr_vec_in_AZ_dqPE7(f_upd_curr_vec_in_AZ_dqPE7) enable((*inhigh*) EN_f_upd_curr_vec_in_AZ_dqPE7) ;
    method f_upd_curr_vec_in_LX_dqPE7(f_upd_curr_vec_in_LX_dqPE7) enable((*inhigh*) EN_f_upd_curr_vec_in_LX_dqPE7) ;
    method f_upd_curr_vec_in_LY_dqPE7(f_upd_curr_vec_in_LY_dqPE7) enable((*inhigh*) EN_f_upd_curr_vec_in_LY_dqPE7) ;
    method f_upd_curr_vec_in_LZ_dqPE7(f_upd_curr_vec_in_LZ_dqPE7) enable((*inhigh*) EN_f_upd_curr_vec_in_LZ_dqPE7) ;
    method dfdq_prev_vec_in_AX_dqPE1(dfdq_prev_vec_in_AX_dqPE1) enable((*inhigh*) EN_dfdq_prev_vec_in_AX_dqPE1) ;
    method dfdq_prev_vec_in_AY_dqPE1(dfdq_prev_vec_in_AY_dqPE1) enable((*inhigh*) EN_dfdq_prev_vec_in_AY_dqPE1) ;
    method dfdq_prev_vec_in_AZ_dqPE1(dfdq_prev_vec_in_AZ_dqPE1) enable((*inhigh*) EN_dfdq_prev_vec_in_AZ_dqPE1) ;
    method dfdq_prev_vec_in_LX_dqPE1(dfdq_prev_vec_in_LX_dqPE1) enable((*inhigh*) EN_dfdq_prev_vec_in_LX_dqPE1) ;
    method dfdq_prev_vec_in_LY_dqPE1(dfdq_prev_vec_in_LY_dqPE1) enable((*inhigh*) EN_dfdq_prev_vec_in_LY_dqPE1) ;
    method dfdq_prev_vec_in_LZ_dqPE1(dfdq_prev_vec_in_LZ_dqPE1) enable((*inhigh*) EN_dfdq_prev_vec_in_LZ_dqPE1) ;
    method dfdq_prev_vec_in_AX_dqPE2(dfdq_prev_vec_in_AX_dqPE2) enable((*inhigh*) EN_dfdq_prev_vec_in_AX_dqPE2) ;
    method dfdq_prev_vec_in_AY_dqPE2(dfdq_prev_vec_in_AY_dqPE2) enable((*inhigh*) EN_dfdq_prev_vec_in_AY_dqPE2) ;
    method dfdq_prev_vec_in_AZ_dqPE2(dfdq_prev_vec_in_AZ_dqPE2) enable((*inhigh*) EN_dfdq_prev_vec_in_AZ_dqPE2) ;
    method dfdq_prev_vec_in_LX_dqPE2(dfdq_prev_vec_in_LX_dqPE2) enable((*inhigh*) EN_dfdq_prev_vec_in_LX_dqPE2) ;
    method dfdq_prev_vec_in_LY_dqPE2(dfdq_prev_vec_in_LY_dqPE2) enable((*inhigh*) EN_dfdq_prev_vec_in_LY_dqPE2) ;
    method dfdq_prev_vec_in_LZ_dqPE2(dfdq_prev_vec_in_LZ_dqPE2) enable((*inhigh*) EN_dfdq_prev_vec_in_LZ_dqPE2) ;
    method dfdq_prev_vec_in_AX_dqPE3(dfdq_prev_vec_in_AX_dqPE3) enable((*inhigh*) EN_dfdq_prev_vec_in_AX_dqPE3) ;
    method dfdq_prev_vec_in_AY_dqPE3(dfdq_prev_vec_in_AY_dqPE3) enable((*inhigh*) EN_dfdq_prev_vec_in_AY_dqPE3) ;
    method dfdq_prev_vec_in_AZ_dqPE3(dfdq_prev_vec_in_AZ_dqPE3) enable((*inhigh*) EN_dfdq_prev_vec_in_AZ_dqPE3) ;
    method dfdq_prev_vec_in_LX_dqPE3(dfdq_prev_vec_in_LX_dqPE3) enable((*inhigh*) EN_dfdq_prev_vec_in_LX_dqPE3) ;
    method dfdq_prev_vec_in_LY_dqPE3(dfdq_prev_vec_in_LY_dqPE3) enable((*inhigh*) EN_dfdq_prev_vec_in_LY_dqPE3) ;
    method dfdq_prev_vec_in_LZ_dqPE3(dfdq_prev_vec_in_LZ_dqPE3) enable((*inhigh*) EN_dfdq_prev_vec_in_LZ_dqPE3) ;
    method dfdq_prev_vec_in_AX_dqPE4(dfdq_prev_vec_in_AX_dqPE4) enable((*inhigh*) EN_dfdq_prev_vec_in_AX_dqPE4) ;
    method dfdq_prev_vec_in_AY_dqPE4(dfdq_prev_vec_in_AY_dqPE4) enable((*inhigh*) EN_dfdq_prev_vec_in_AY_dqPE4) ;
    method dfdq_prev_vec_in_AZ_dqPE4(dfdq_prev_vec_in_AZ_dqPE4) enable((*inhigh*) EN_dfdq_prev_vec_in_AZ_dqPE4) ;
    method dfdq_prev_vec_in_LX_dqPE4(dfdq_prev_vec_in_LX_dqPE4) enable((*inhigh*) EN_dfdq_prev_vec_in_LX_dqPE4) ;
    method dfdq_prev_vec_in_LY_dqPE4(dfdq_prev_vec_in_LY_dqPE4) enable((*inhigh*) EN_dfdq_prev_vec_in_LY_dqPE4) ;
    method dfdq_prev_vec_in_LZ_dqPE4(dfdq_prev_vec_in_LZ_dqPE4) enable((*inhigh*) EN_dfdq_prev_vec_in_LZ_dqPE4) ;
    method dfdq_prev_vec_in_AX_dqPE5(dfdq_prev_vec_in_AX_dqPE5) enable((*inhigh*) EN_dfdq_prev_vec_in_AX_dqPE5) ;
    method dfdq_prev_vec_in_AY_dqPE5(dfdq_prev_vec_in_AY_dqPE5) enable((*inhigh*) EN_dfdq_prev_vec_in_AY_dqPE5) ;
    method dfdq_prev_vec_in_AZ_dqPE5(dfdq_prev_vec_in_AZ_dqPE5) enable((*inhigh*) EN_dfdq_prev_vec_in_AZ_dqPE5) ;
    method dfdq_prev_vec_in_LX_dqPE5(dfdq_prev_vec_in_LX_dqPE5) enable((*inhigh*) EN_dfdq_prev_vec_in_LX_dqPE5) ;
    method dfdq_prev_vec_in_LY_dqPE5(dfdq_prev_vec_in_LY_dqPE5) enable((*inhigh*) EN_dfdq_prev_vec_in_LY_dqPE5) ;
    method dfdq_prev_vec_in_LZ_dqPE5(dfdq_prev_vec_in_LZ_dqPE5) enable((*inhigh*) EN_dfdq_prev_vec_in_LZ_dqPE5) ;
    method dfdq_prev_vec_in_AX_dqPE6(dfdq_prev_vec_in_AX_dqPE6) enable((*inhigh*) EN_dfdq_prev_vec_in_AX_dqPE6) ;
    method dfdq_prev_vec_in_AY_dqPE6(dfdq_prev_vec_in_AY_dqPE6) enable((*inhigh*) EN_dfdq_prev_vec_in_AY_dqPE6) ;
    method dfdq_prev_vec_in_AZ_dqPE6(dfdq_prev_vec_in_AZ_dqPE6) enable((*inhigh*) EN_dfdq_prev_vec_in_AZ_dqPE6) ;
    method dfdq_prev_vec_in_LX_dqPE6(dfdq_prev_vec_in_LX_dqPE6) enable((*inhigh*) EN_dfdq_prev_vec_in_LX_dqPE6) ;
    method dfdq_prev_vec_in_LY_dqPE6(dfdq_prev_vec_in_LY_dqPE6) enable((*inhigh*) EN_dfdq_prev_vec_in_LY_dqPE6) ;
    method dfdq_prev_vec_in_LZ_dqPE6(dfdq_prev_vec_in_LZ_dqPE6) enable((*inhigh*) EN_dfdq_prev_vec_in_LZ_dqPE6) ;
    method dfdq_prev_vec_in_AX_dqPE7(dfdq_prev_vec_in_AX_dqPE7) enable((*inhigh*) EN_dfdq_prev_vec_in_AX_dqPE7) ;
    method dfdq_prev_vec_in_AY_dqPE7(dfdq_prev_vec_in_AY_dqPE7) enable((*inhigh*) EN_dfdq_prev_vec_in_AY_dqPE7) ;
    method dfdq_prev_vec_in_AZ_dqPE7(dfdq_prev_vec_in_AZ_dqPE7) enable((*inhigh*) EN_dfdq_prev_vec_in_AZ_dqPE7) ;
    method dfdq_prev_vec_in_LX_dqPE7(dfdq_prev_vec_in_LX_dqPE7) enable((*inhigh*) EN_dfdq_prev_vec_in_LX_dqPE7) ;
    method dfdq_prev_vec_in_LY_dqPE7(dfdq_prev_vec_in_LY_dqPE7) enable((*inhigh*) EN_dfdq_prev_vec_in_LY_dqPE7) ;
    method dfdq_prev_vec_in_LZ_dqPE7(dfdq_prev_vec_in_LZ_dqPE7) enable((*inhigh*) EN_dfdq_prev_vec_in_LZ_dqPE7) ;
    method dfdq_upd_curr_vec_in_AX_dqPE1(dfdq_upd_curr_vec_in_AX_dqPE1) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AX_dqPE1) ;
    method dfdq_upd_curr_vec_in_AY_dqPE1(dfdq_upd_curr_vec_in_AY_dqPE1) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AY_dqPE1) ;
    method dfdq_upd_curr_vec_in_AZ_dqPE1(dfdq_upd_curr_vec_in_AZ_dqPE1) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AZ_dqPE1) ;
    method dfdq_upd_curr_vec_in_LX_dqPE1(dfdq_upd_curr_vec_in_LX_dqPE1) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LX_dqPE1) ;
    method dfdq_upd_curr_vec_in_LY_dqPE1(dfdq_upd_curr_vec_in_LY_dqPE1) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LY_dqPE1) ;
    method dfdq_upd_curr_vec_in_LZ_dqPE1(dfdq_upd_curr_vec_in_LZ_dqPE1) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LZ_dqPE1) ;
    method dfdq_upd_curr_vec_in_AX_dqPE2(dfdq_upd_curr_vec_in_AX_dqPE2) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AX_dqPE2) ;
    method dfdq_upd_curr_vec_in_AY_dqPE2(dfdq_upd_curr_vec_in_AY_dqPE2) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AY_dqPE2) ;
    method dfdq_upd_curr_vec_in_AZ_dqPE2(dfdq_upd_curr_vec_in_AZ_dqPE2) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AZ_dqPE2) ;
    method dfdq_upd_curr_vec_in_LX_dqPE2(dfdq_upd_curr_vec_in_LX_dqPE2) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LX_dqPE2) ;
    method dfdq_upd_curr_vec_in_LY_dqPE2(dfdq_upd_curr_vec_in_LY_dqPE2) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LY_dqPE2) ;
    method dfdq_upd_curr_vec_in_LZ_dqPE2(dfdq_upd_curr_vec_in_LZ_dqPE2) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LZ_dqPE2) ;
    method dfdq_upd_curr_vec_in_AX_dqPE3(dfdq_upd_curr_vec_in_AX_dqPE3) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AX_dqPE3) ;
    method dfdq_upd_curr_vec_in_AY_dqPE3(dfdq_upd_curr_vec_in_AY_dqPE3) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AY_dqPE3) ;
    method dfdq_upd_curr_vec_in_AZ_dqPE3(dfdq_upd_curr_vec_in_AZ_dqPE3) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AZ_dqPE3) ;
    method dfdq_upd_curr_vec_in_LX_dqPE3(dfdq_upd_curr_vec_in_LX_dqPE3) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LX_dqPE3) ;
    method dfdq_upd_curr_vec_in_LY_dqPE3(dfdq_upd_curr_vec_in_LY_dqPE3) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LY_dqPE3) ;
    method dfdq_upd_curr_vec_in_LZ_dqPE3(dfdq_upd_curr_vec_in_LZ_dqPE3) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LZ_dqPE3) ;
    method dfdq_upd_curr_vec_in_AX_dqPE4(dfdq_upd_curr_vec_in_AX_dqPE4) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AX_dqPE4) ;
    method dfdq_upd_curr_vec_in_AY_dqPE4(dfdq_upd_curr_vec_in_AY_dqPE4) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AY_dqPE4) ;
    method dfdq_upd_curr_vec_in_AZ_dqPE4(dfdq_upd_curr_vec_in_AZ_dqPE4) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AZ_dqPE4) ;
    method dfdq_upd_curr_vec_in_LX_dqPE4(dfdq_upd_curr_vec_in_LX_dqPE4) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LX_dqPE4) ;
    method dfdq_upd_curr_vec_in_LY_dqPE4(dfdq_upd_curr_vec_in_LY_dqPE4) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LY_dqPE4) ;
    method dfdq_upd_curr_vec_in_LZ_dqPE4(dfdq_upd_curr_vec_in_LZ_dqPE4) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LZ_dqPE4) ;
    method dfdq_upd_curr_vec_in_AX_dqPE5(dfdq_upd_curr_vec_in_AX_dqPE5) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AX_dqPE5) ;
    method dfdq_upd_curr_vec_in_AY_dqPE5(dfdq_upd_curr_vec_in_AY_dqPE5) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AY_dqPE5) ;
    method dfdq_upd_curr_vec_in_AZ_dqPE5(dfdq_upd_curr_vec_in_AZ_dqPE5) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AZ_dqPE5) ;
    method dfdq_upd_curr_vec_in_LX_dqPE5(dfdq_upd_curr_vec_in_LX_dqPE5) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LX_dqPE5) ;
    method dfdq_upd_curr_vec_in_LY_dqPE5(dfdq_upd_curr_vec_in_LY_dqPE5) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LY_dqPE5) ;
    method dfdq_upd_curr_vec_in_LZ_dqPE5(dfdq_upd_curr_vec_in_LZ_dqPE5) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LZ_dqPE5) ;
    method dfdq_upd_curr_vec_in_AX_dqPE6(dfdq_upd_curr_vec_in_AX_dqPE6) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AX_dqPE6) ;
    method dfdq_upd_curr_vec_in_AY_dqPE6(dfdq_upd_curr_vec_in_AY_dqPE6) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AY_dqPE6) ;
    method dfdq_upd_curr_vec_in_AZ_dqPE6(dfdq_upd_curr_vec_in_AZ_dqPE6) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AZ_dqPE6) ;
    method dfdq_upd_curr_vec_in_LX_dqPE6(dfdq_upd_curr_vec_in_LX_dqPE6) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LX_dqPE6) ;
    method dfdq_upd_curr_vec_in_LY_dqPE6(dfdq_upd_curr_vec_in_LY_dqPE6) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LY_dqPE6) ;
    method dfdq_upd_curr_vec_in_LZ_dqPE6(dfdq_upd_curr_vec_in_LZ_dqPE6) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LZ_dqPE6) ;
    method dfdq_upd_curr_vec_in_AX_dqPE7(dfdq_upd_curr_vec_in_AX_dqPE7) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AX_dqPE7) ;
    method dfdq_upd_curr_vec_in_AY_dqPE7(dfdq_upd_curr_vec_in_AY_dqPE7) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AY_dqPE7) ;
    method dfdq_upd_curr_vec_in_AZ_dqPE7(dfdq_upd_curr_vec_in_AZ_dqPE7) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_AZ_dqPE7) ;
    method dfdq_upd_curr_vec_in_LX_dqPE7(dfdq_upd_curr_vec_in_LX_dqPE7) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LX_dqPE7) ;
    method dfdq_upd_curr_vec_in_LY_dqPE7(dfdq_upd_curr_vec_in_LY_dqPE7) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LY_dqPE7) ;
    method dfdq_upd_curr_vec_in_LZ_dqPE7(dfdq_upd_curr_vec_in_LZ_dqPE7) enable((*inhigh*) EN_dfdq_upd_curr_vec_in_LZ_dqPE7) ;
    method dfdqd_prev_vec_in_AX_dqdPE1(dfdqd_prev_vec_in_AX_dqdPE1) enable((*inhigh*) EN_dfdqd_prev_vec_in_AX_dqdPE1) ;
    method dfdqd_prev_vec_in_AY_dqdPE1(dfdqd_prev_vec_in_AY_dqdPE1) enable((*inhigh*) EN_dfdqd_prev_vec_in_AY_dqdPE1) ;
    method dfdqd_prev_vec_in_AZ_dqdPE1(dfdqd_prev_vec_in_AZ_dqdPE1) enable((*inhigh*) EN_dfdqd_prev_vec_in_AZ_dqdPE1) ;
    method dfdqd_prev_vec_in_LX_dqdPE1(dfdqd_prev_vec_in_LX_dqdPE1) enable((*inhigh*) EN_dfdqd_prev_vec_in_LX_dqdPE1) ;
    method dfdqd_prev_vec_in_LY_dqdPE1(dfdqd_prev_vec_in_LY_dqdPE1) enable((*inhigh*) EN_dfdqd_prev_vec_in_LY_dqdPE1) ;
    method dfdqd_prev_vec_in_LZ_dqdPE1(dfdqd_prev_vec_in_LZ_dqdPE1) enable((*inhigh*) EN_dfdqd_prev_vec_in_LZ_dqdPE1) ;
    method dfdqd_prev_vec_in_AX_dqdPE2(dfdqd_prev_vec_in_AX_dqdPE2) enable((*inhigh*) EN_dfdqd_prev_vec_in_AX_dqdPE2) ;
    method dfdqd_prev_vec_in_AY_dqdPE2(dfdqd_prev_vec_in_AY_dqdPE2) enable((*inhigh*) EN_dfdqd_prev_vec_in_AY_dqdPE2) ;
    method dfdqd_prev_vec_in_AZ_dqdPE2(dfdqd_prev_vec_in_AZ_dqdPE2) enable((*inhigh*) EN_dfdqd_prev_vec_in_AZ_dqdPE2) ;
    method dfdqd_prev_vec_in_LX_dqdPE2(dfdqd_prev_vec_in_LX_dqdPE2) enable((*inhigh*) EN_dfdqd_prev_vec_in_LX_dqdPE2) ;
    method dfdqd_prev_vec_in_LY_dqdPE2(dfdqd_prev_vec_in_LY_dqdPE2) enable((*inhigh*) EN_dfdqd_prev_vec_in_LY_dqdPE2) ;
    method dfdqd_prev_vec_in_LZ_dqdPE2(dfdqd_prev_vec_in_LZ_dqdPE2) enable((*inhigh*) EN_dfdqd_prev_vec_in_LZ_dqdPE2) ;
    method dfdqd_prev_vec_in_AX_dqdPE3(dfdqd_prev_vec_in_AX_dqdPE3) enable((*inhigh*) EN_dfdqd_prev_vec_in_AX_dqdPE3) ;
    method dfdqd_prev_vec_in_AY_dqdPE3(dfdqd_prev_vec_in_AY_dqdPE3) enable((*inhigh*) EN_dfdqd_prev_vec_in_AY_dqdPE3) ;
    method dfdqd_prev_vec_in_AZ_dqdPE3(dfdqd_prev_vec_in_AZ_dqdPE3) enable((*inhigh*) EN_dfdqd_prev_vec_in_AZ_dqdPE3) ;
    method dfdqd_prev_vec_in_LX_dqdPE3(dfdqd_prev_vec_in_LX_dqdPE3) enable((*inhigh*) EN_dfdqd_prev_vec_in_LX_dqdPE3) ;
    method dfdqd_prev_vec_in_LY_dqdPE3(dfdqd_prev_vec_in_LY_dqdPE3) enable((*inhigh*) EN_dfdqd_prev_vec_in_LY_dqdPE3) ;
    method dfdqd_prev_vec_in_LZ_dqdPE3(dfdqd_prev_vec_in_LZ_dqdPE3) enable((*inhigh*) EN_dfdqd_prev_vec_in_LZ_dqdPE3) ;
    method dfdqd_prev_vec_in_AX_dqdPE4(dfdqd_prev_vec_in_AX_dqdPE4) enable((*inhigh*) EN_dfdqd_prev_vec_in_AX_dqdPE4) ;
    method dfdqd_prev_vec_in_AY_dqdPE4(dfdqd_prev_vec_in_AY_dqdPE4) enable((*inhigh*) EN_dfdqd_prev_vec_in_AY_dqdPE4) ;
    method dfdqd_prev_vec_in_AZ_dqdPE4(dfdqd_prev_vec_in_AZ_dqdPE4) enable((*inhigh*) EN_dfdqd_prev_vec_in_AZ_dqdPE4) ;
    method dfdqd_prev_vec_in_LX_dqdPE4(dfdqd_prev_vec_in_LX_dqdPE4) enable((*inhigh*) EN_dfdqd_prev_vec_in_LX_dqdPE4) ;
    method dfdqd_prev_vec_in_LY_dqdPE4(dfdqd_prev_vec_in_LY_dqdPE4) enable((*inhigh*) EN_dfdqd_prev_vec_in_LY_dqdPE4) ;
    method dfdqd_prev_vec_in_LZ_dqdPE4(dfdqd_prev_vec_in_LZ_dqdPE4) enable((*inhigh*) EN_dfdqd_prev_vec_in_LZ_dqdPE4) ;
    method dfdqd_prev_vec_in_AX_dqdPE5(dfdqd_prev_vec_in_AX_dqdPE5) enable((*inhigh*) EN_dfdqd_prev_vec_in_AX_dqdPE5) ;
    method dfdqd_prev_vec_in_AY_dqdPE5(dfdqd_prev_vec_in_AY_dqdPE5) enable((*inhigh*) EN_dfdqd_prev_vec_in_AY_dqdPE5) ;
    method dfdqd_prev_vec_in_AZ_dqdPE5(dfdqd_prev_vec_in_AZ_dqdPE5) enable((*inhigh*) EN_dfdqd_prev_vec_in_AZ_dqdPE5) ;
    method dfdqd_prev_vec_in_LX_dqdPE5(dfdqd_prev_vec_in_LX_dqdPE5) enable((*inhigh*) EN_dfdqd_prev_vec_in_LX_dqdPE5) ;
    method dfdqd_prev_vec_in_LY_dqdPE5(dfdqd_prev_vec_in_LY_dqdPE5) enable((*inhigh*) EN_dfdqd_prev_vec_in_LY_dqdPE5) ;
    method dfdqd_prev_vec_in_LZ_dqdPE5(dfdqd_prev_vec_in_LZ_dqdPE5) enable((*inhigh*) EN_dfdqd_prev_vec_in_LZ_dqdPE5) ;
    method dfdqd_prev_vec_in_AX_dqdPE6(dfdqd_prev_vec_in_AX_dqdPE6) enable((*inhigh*) EN_dfdqd_prev_vec_in_AX_dqdPE6) ;
    method dfdqd_prev_vec_in_AY_dqdPE6(dfdqd_prev_vec_in_AY_dqdPE6) enable((*inhigh*) EN_dfdqd_prev_vec_in_AY_dqdPE6) ;
    method dfdqd_prev_vec_in_AZ_dqdPE6(dfdqd_prev_vec_in_AZ_dqdPE6) enable((*inhigh*) EN_dfdqd_prev_vec_in_AZ_dqdPE6) ;
    method dfdqd_prev_vec_in_LX_dqdPE6(dfdqd_prev_vec_in_LX_dqdPE6) enable((*inhigh*) EN_dfdqd_prev_vec_in_LX_dqdPE6) ;
    method dfdqd_prev_vec_in_LY_dqdPE6(dfdqd_prev_vec_in_LY_dqdPE6) enable((*inhigh*) EN_dfdqd_prev_vec_in_LY_dqdPE6) ;
    method dfdqd_prev_vec_in_LZ_dqdPE6(dfdqd_prev_vec_in_LZ_dqdPE6) enable((*inhigh*) EN_dfdqd_prev_vec_in_LZ_dqdPE6) ;
    method dfdqd_prev_vec_in_AX_dqdPE7(dfdqd_prev_vec_in_AX_dqdPE7) enable((*inhigh*) EN_dfdqd_prev_vec_in_AX_dqdPE7) ;
    method dfdqd_prev_vec_in_AY_dqdPE7(dfdqd_prev_vec_in_AY_dqdPE7) enable((*inhigh*) EN_dfdqd_prev_vec_in_AY_dqdPE7) ;
    method dfdqd_prev_vec_in_AZ_dqdPE7(dfdqd_prev_vec_in_AZ_dqdPE7) enable((*inhigh*) EN_dfdqd_prev_vec_in_AZ_dqdPE7) ;
    method dfdqd_prev_vec_in_LX_dqdPE7(dfdqd_prev_vec_in_LX_dqdPE7) enable((*inhigh*) EN_dfdqd_prev_vec_in_LX_dqdPE7) ;
    method dfdqd_prev_vec_in_LY_dqdPE7(dfdqd_prev_vec_in_LY_dqdPE7) enable((*inhigh*) EN_dfdqd_prev_vec_in_LY_dqdPE7) ;
    method dfdqd_prev_vec_in_LZ_dqdPE7(dfdqd_prev_vec_in_LZ_dqdPE7) enable((*inhigh*) EN_dfdqd_prev_vec_in_LZ_dqdPE7) ;
    method dfdqd_upd_curr_vec_in_AX_dqdPE1(dfdqd_upd_curr_vec_in_AX_dqdPE1) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AX_dqdPE1) ;
    method dfdqd_upd_curr_vec_in_AY_dqdPE1(dfdqd_upd_curr_vec_in_AY_dqdPE1) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AY_dqdPE1) ;
    method dfdqd_upd_curr_vec_in_AZ_dqdPE1(dfdqd_upd_curr_vec_in_AZ_dqdPE1) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AZ_dqdPE1) ;
    method dfdqd_upd_curr_vec_in_LX_dqdPE1(dfdqd_upd_curr_vec_in_LX_dqdPE1) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LX_dqdPE1) ;
    method dfdqd_upd_curr_vec_in_LY_dqdPE1(dfdqd_upd_curr_vec_in_LY_dqdPE1) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LY_dqdPE1) ;
    method dfdqd_upd_curr_vec_in_LZ_dqdPE1(dfdqd_upd_curr_vec_in_LZ_dqdPE1) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LZ_dqdPE1) ;
    method dfdqd_upd_curr_vec_in_AX_dqdPE2(dfdqd_upd_curr_vec_in_AX_dqdPE2) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AX_dqdPE2) ;
    method dfdqd_upd_curr_vec_in_AY_dqdPE2(dfdqd_upd_curr_vec_in_AY_dqdPE2) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AY_dqdPE2) ;
    method dfdqd_upd_curr_vec_in_AZ_dqdPE2(dfdqd_upd_curr_vec_in_AZ_dqdPE2) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AZ_dqdPE2) ;
    method dfdqd_upd_curr_vec_in_LX_dqdPE2(dfdqd_upd_curr_vec_in_LX_dqdPE2) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LX_dqdPE2) ;
    method dfdqd_upd_curr_vec_in_LY_dqdPE2(dfdqd_upd_curr_vec_in_LY_dqdPE2) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LY_dqdPE2) ;
    method dfdqd_upd_curr_vec_in_LZ_dqdPE2(dfdqd_upd_curr_vec_in_LZ_dqdPE2) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LZ_dqdPE2) ;
    method dfdqd_upd_curr_vec_in_AX_dqdPE3(dfdqd_upd_curr_vec_in_AX_dqdPE3) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AX_dqdPE3) ;
    method dfdqd_upd_curr_vec_in_AY_dqdPE3(dfdqd_upd_curr_vec_in_AY_dqdPE3) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AY_dqdPE3) ;
    method dfdqd_upd_curr_vec_in_AZ_dqdPE3(dfdqd_upd_curr_vec_in_AZ_dqdPE3) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AZ_dqdPE3) ;
    method dfdqd_upd_curr_vec_in_LX_dqdPE3(dfdqd_upd_curr_vec_in_LX_dqdPE3) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LX_dqdPE3) ;
    method dfdqd_upd_curr_vec_in_LY_dqdPE3(dfdqd_upd_curr_vec_in_LY_dqdPE3) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LY_dqdPE3) ;
    method dfdqd_upd_curr_vec_in_LZ_dqdPE3(dfdqd_upd_curr_vec_in_LZ_dqdPE3) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LZ_dqdPE3) ;
    method dfdqd_upd_curr_vec_in_AX_dqdPE4(dfdqd_upd_curr_vec_in_AX_dqdPE4) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AX_dqdPE4) ;
    method dfdqd_upd_curr_vec_in_AY_dqdPE4(dfdqd_upd_curr_vec_in_AY_dqdPE4) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AY_dqdPE4) ;
    method dfdqd_upd_curr_vec_in_AZ_dqdPE4(dfdqd_upd_curr_vec_in_AZ_dqdPE4) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AZ_dqdPE4) ;
    method dfdqd_upd_curr_vec_in_LX_dqdPE4(dfdqd_upd_curr_vec_in_LX_dqdPE4) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LX_dqdPE4) ;
    method dfdqd_upd_curr_vec_in_LY_dqdPE4(dfdqd_upd_curr_vec_in_LY_dqdPE4) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LY_dqdPE4) ;
    method dfdqd_upd_curr_vec_in_LZ_dqdPE4(dfdqd_upd_curr_vec_in_LZ_dqdPE4) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LZ_dqdPE4) ;
    method dfdqd_upd_curr_vec_in_AX_dqdPE5(dfdqd_upd_curr_vec_in_AX_dqdPE5) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AX_dqdPE5) ;
    method dfdqd_upd_curr_vec_in_AY_dqdPE5(dfdqd_upd_curr_vec_in_AY_dqdPE5) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AY_dqdPE5) ;
    method dfdqd_upd_curr_vec_in_AZ_dqdPE5(dfdqd_upd_curr_vec_in_AZ_dqdPE5) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AZ_dqdPE5) ;
    method dfdqd_upd_curr_vec_in_LX_dqdPE5(dfdqd_upd_curr_vec_in_LX_dqdPE5) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LX_dqdPE5) ;
    method dfdqd_upd_curr_vec_in_LY_dqdPE5(dfdqd_upd_curr_vec_in_LY_dqdPE5) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LY_dqdPE5) ;
    method dfdqd_upd_curr_vec_in_LZ_dqdPE5(dfdqd_upd_curr_vec_in_LZ_dqdPE5) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LZ_dqdPE5) ;
    method dfdqd_upd_curr_vec_in_AX_dqdPE6(dfdqd_upd_curr_vec_in_AX_dqdPE6) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AX_dqdPE6) ;
    method dfdqd_upd_curr_vec_in_AY_dqdPE6(dfdqd_upd_curr_vec_in_AY_dqdPE6) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AY_dqdPE6) ;
    method dfdqd_upd_curr_vec_in_AZ_dqdPE6(dfdqd_upd_curr_vec_in_AZ_dqdPE6) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AZ_dqdPE6) ;
    method dfdqd_upd_curr_vec_in_LX_dqdPE6(dfdqd_upd_curr_vec_in_LX_dqdPE6) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LX_dqdPE6) ;
    method dfdqd_upd_curr_vec_in_LY_dqdPE6(dfdqd_upd_curr_vec_in_LY_dqdPE6) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LY_dqdPE6) ;
    method dfdqd_upd_curr_vec_in_LZ_dqdPE6(dfdqd_upd_curr_vec_in_LZ_dqdPE6) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LZ_dqdPE6) ;
    method dfdqd_upd_curr_vec_in_AX_dqdPE7(dfdqd_upd_curr_vec_in_AX_dqdPE7) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AX_dqdPE7) ;
    method dfdqd_upd_curr_vec_in_AY_dqdPE7(dfdqd_upd_curr_vec_in_AY_dqdPE7) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AY_dqdPE7) ;
    method dfdqd_upd_curr_vec_in_AZ_dqdPE7(dfdqd_upd_curr_vec_in_AZ_dqdPE7) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_AZ_dqdPE7) ;
    method dfdqd_upd_curr_vec_in_LX_dqdPE7(dfdqd_upd_curr_vec_in_LX_dqdPE7) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LX_dqdPE7) ;
    method dfdqd_upd_curr_vec_in_LY_dqdPE7(dfdqd_upd_curr_vec_in_LY_dqdPE7) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LY_dqdPE7) ;
    method dfdqd_upd_curr_vec_in_LZ_dqdPE7(dfdqd_upd_curr_vec_in_LZ_dqdPE7) enable((*inhigh*) EN_dfdqd_upd_curr_vec_in_LZ_dqdPE7) ;

    method minv_block_in_R1_C1_dqdPE1(minv_block_in_R1_C1_dqdPE1) enable((*inhigh*) EN_minv_block_in_R1_C1_dqdPE1) ;
    method minv_block_in_R2_C1_dqdPE1(minv_block_in_R2_C1_dqdPE1) enable((*inhigh*) EN_minv_block_in_R2_C1_dqdPE1) ;
    method minv_block_in_R3_C1_dqdPE1(minv_block_in_R3_C1_dqdPE1) enable((*inhigh*) EN_minv_block_in_R3_C1_dqdPE1) ;
    method minv_block_in_R4_C1_dqdPE1(minv_block_in_R4_C1_dqdPE1) enable((*inhigh*) EN_minv_block_in_R4_C1_dqdPE1) ;
    method minv_block_in_R5_C1_dqdPE1(minv_block_in_R5_C1_dqdPE1) enable((*inhigh*) EN_minv_block_in_R5_C1_dqdPE1) ;
    method minv_block_in_R6_C1_dqdPE1(minv_block_in_R6_C1_dqdPE1) enable((*inhigh*) EN_minv_block_in_R6_C1_dqdPE1) ;
    method minv_block_in_R7_C1_dqdPE1(minv_block_in_R7_C1_dqdPE1) enable((*inhigh*) EN_minv_block_in_R7_C1_dqdPE1) ;
    method minv_block_in_R1_C2_dqdPE1(minv_block_in_R1_C2_dqdPE1) enable((*inhigh*) EN_minv_block_in_R1_C2_dqdPE1) ;
    method minv_block_in_R2_C2_dqdPE1(minv_block_in_R2_C2_dqdPE1) enable((*inhigh*) EN_minv_block_in_R2_C2_dqdPE1) ;
    method minv_block_in_R3_C2_dqdPE1(minv_block_in_R3_C2_dqdPE1) enable((*inhigh*) EN_minv_block_in_R3_C2_dqdPE1) ;
    method minv_block_in_R4_C2_dqdPE1(minv_block_in_R4_C2_dqdPE1) enable((*inhigh*) EN_minv_block_in_R4_C2_dqdPE1) ;
    method minv_block_in_R5_C2_dqdPE1(minv_block_in_R5_C2_dqdPE1) enable((*inhigh*) EN_minv_block_in_R5_C2_dqdPE1) ;
    method minv_block_in_R6_C2_dqdPE1(minv_block_in_R6_C2_dqdPE1) enable((*inhigh*) EN_minv_block_in_R6_C2_dqdPE1) ;
    method minv_block_in_R7_C2_dqdPE1(minv_block_in_R7_C2_dqdPE1) enable((*inhigh*) EN_minv_block_in_R7_C2_dqdPE1) ;
    method minv_block_in_R1_C3_dqdPE1(minv_block_in_R1_C3_dqdPE1) enable((*inhigh*) EN_minv_block_in_R1_C3_dqdPE1) ;
    method minv_block_in_R2_C3_dqdPE1(minv_block_in_R2_C3_dqdPE1) enable((*inhigh*) EN_minv_block_in_R2_C3_dqdPE1) ;
    method minv_block_in_R3_C3_dqdPE1(minv_block_in_R3_C3_dqdPE1) enable((*inhigh*) EN_minv_block_in_R3_C3_dqdPE1) ;
    method minv_block_in_R4_C3_dqdPE1(minv_block_in_R4_C3_dqdPE1) enable((*inhigh*) EN_minv_block_in_R4_C3_dqdPE1) ;
    method minv_block_in_R5_C3_dqdPE1(minv_block_in_R5_C3_dqdPE1) enable((*inhigh*) EN_minv_block_in_R5_C3_dqdPE1) ;
    method minv_block_in_R6_C3_dqdPE1(minv_block_in_R6_C3_dqdPE1) enable((*inhigh*) EN_minv_block_in_R6_C3_dqdPE1) ;
    method minv_block_in_R7_C3_dqdPE1(minv_block_in_R7_C3_dqdPE1) enable((*inhigh*) EN_minv_block_in_R7_C3_dqdPE1) ;
    method minv_block_in_R1_C4_dqdPE1(minv_block_in_R1_C4_dqdPE1) enable((*inhigh*) EN_minv_block_in_R1_C4_dqdPE1) ;
    method minv_block_in_R2_C4_dqdPE1(minv_block_in_R2_C4_dqdPE1) enable((*inhigh*) EN_minv_block_in_R2_C4_dqdPE1) ;
    method minv_block_in_R3_C4_dqdPE1(minv_block_in_R3_C4_dqdPE1) enable((*inhigh*) EN_minv_block_in_R3_C4_dqdPE1) ;
    method minv_block_in_R4_C4_dqdPE1(minv_block_in_R4_C4_dqdPE1) enable((*inhigh*) EN_minv_block_in_R4_C4_dqdPE1) ;
    method minv_block_in_R5_C4_dqdPE1(minv_block_in_R5_C4_dqdPE1) enable((*inhigh*) EN_minv_block_in_R5_C4_dqdPE1) ;
    method minv_block_in_R6_C4_dqdPE1(minv_block_in_R6_C4_dqdPE1) enable((*inhigh*) EN_minv_block_in_R6_C4_dqdPE1) ;
    method minv_block_in_R7_C4_dqdPE1(minv_block_in_R7_C4_dqdPE1) enable((*inhigh*) EN_minv_block_in_R7_C4_dqdPE1) ;
    method minv_block_in_R1_C5_dqdPE1(minv_block_in_R1_C5_dqdPE1) enable((*inhigh*) EN_minv_block_in_R1_C5_dqdPE1) ;
    method minv_block_in_R2_C5_dqdPE1(minv_block_in_R2_C5_dqdPE1) enable((*inhigh*) EN_minv_block_in_R2_C5_dqdPE1) ;
    method minv_block_in_R3_C5_dqdPE1(minv_block_in_R3_C5_dqdPE1) enable((*inhigh*) EN_minv_block_in_R3_C5_dqdPE1) ;
    method minv_block_in_R4_C5_dqdPE1(minv_block_in_R4_C5_dqdPE1) enable((*inhigh*) EN_minv_block_in_R4_C5_dqdPE1) ;
    method minv_block_in_R5_C5_dqdPE1(minv_block_in_R5_C5_dqdPE1) enable((*inhigh*) EN_minv_block_in_R5_C5_dqdPE1) ;
    method minv_block_in_R6_C5_dqdPE1(minv_block_in_R6_C5_dqdPE1) enable((*inhigh*) EN_minv_block_in_R6_C5_dqdPE1) ;
    method minv_block_in_R7_C5_dqdPE1(minv_block_in_R7_C5_dqdPE1) enable((*inhigh*) EN_minv_block_in_R7_C5_dqdPE1) ;
    method minv_block_in_R1_C6_dqdPE1(minv_block_in_R1_C6_dqdPE1) enable((*inhigh*) EN_minv_block_in_R1_C6_dqdPE1) ;
    method minv_block_in_R2_C6_dqdPE1(minv_block_in_R2_C6_dqdPE1) enable((*inhigh*) EN_minv_block_in_R2_C6_dqdPE1) ;
    method minv_block_in_R3_C6_dqdPE1(minv_block_in_R3_C6_dqdPE1) enable((*inhigh*) EN_minv_block_in_R3_C6_dqdPE1) ;
    method minv_block_in_R4_C6_dqdPE1(minv_block_in_R4_C6_dqdPE1) enable((*inhigh*) EN_minv_block_in_R4_C6_dqdPE1) ;
    method minv_block_in_R5_C6_dqdPE1(minv_block_in_R5_C6_dqdPE1) enable((*inhigh*) EN_minv_block_in_R5_C6_dqdPE1) ;
    method minv_block_in_R6_C6_dqdPE1(minv_block_in_R6_C6_dqdPE1) enable((*inhigh*) EN_minv_block_in_R6_C6_dqdPE1) ;
    method minv_block_in_R7_C6_dqdPE1(minv_block_in_R7_C6_dqdPE1) enable((*inhigh*) EN_minv_block_in_R7_C6_dqdPE1) ;
    method minv_block_in_R1_C7_dqdPE1(minv_block_in_R1_C7_dqdPE1) enable((*inhigh*) EN_minv_block_in_R1_C7_dqdPE1) ;
    method minv_block_in_R2_C7_dqdPE1(minv_block_in_R2_C7_dqdPE1) enable((*inhigh*) EN_minv_block_in_R2_C7_dqdPE1) ;
    method minv_block_in_R3_C7_dqdPE1(minv_block_in_R3_C7_dqdPE1) enable((*inhigh*) EN_minv_block_in_R3_C7_dqdPE1) ;
    method minv_block_in_R4_C7_dqdPE1(minv_block_in_R4_C7_dqdPE1) enable((*inhigh*) EN_minv_block_in_R4_C7_dqdPE1) ;
    method minv_block_in_R5_C7_dqdPE1(minv_block_in_R5_C7_dqdPE1) enable((*inhigh*) EN_minv_block_in_R5_C7_dqdPE1) ;
    method minv_block_in_R6_C7_dqdPE1(minv_block_in_R6_C7_dqdPE1) enable((*inhigh*) EN_minv_block_in_R6_C7_dqdPE1) ;
    method minv_block_in_R7_C7_dqdPE1(minv_block_in_R7_C7_dqdPE1) enable((*inhigh*) EN_minv_block_in_R7_C7_dqdPE1) ;
    method minv_block_in_R1_C1_dqdPE2(minv_block_in_R1_C1_dqdPE2) enable((*inhigh*) EN_minv_block_in_R1_C1_dqdPE2) ;
    method minv_block_in_R2_C1_dqdPE2(minv_block_in_R2_C1_dqdPE2) enable((*inhigh*) EN_minv_block_in_R2_C1_dqdPE2) ;
    method minv_block_in_R3_C1_dqdPE2(minv_block_in_R3_C1_dqdPE2) enable((*inhigh*) EN_minv_block_in_R3_C1_dqdPE2) ;
    method minv_block_in_R4_C1_dqdPE2(minv_block_in_R4_C1_dqdPE2) enable((*inhigh*) EN_minv_block_in_R4_C1_dqdPE2) ;
    method minv_block_in_R5_C1_dqdPE2(minv_block_in_R5_C1_dqdPE2) enable((*inhigh*) EN_minv_block_in_R5_C1_dqdPE2) ;
    method minv_block_in_R6_C1_dqdPE2(minv_block_in_R6_C1_dqdPE2) enable((*inhigh*) EN_minv_block_in_R6_C1_dqdPE2) ;
    method minv_block_in_R7_C1_dqdPE2(minv_block_in_R7_C1_dqdPE2) enable((*inhigh*) EN_minv_block_in_R7_C1_dqdPE2) ;
    method minv_block_in_R1_C2_dqdPE2(minv_block_in_R1_C2_dqdPE2) enable((*inhigh*) EN_minv_block_in_R1_C2_dqdPE2) ;
    method minv_block_in_R2_C2_dqdPE2(minv_block_in_R2_C2_dqdPE2) enable((*inhigh*) EN_minv_block_in_R2_C2_dqdPE2) ;
    method minv_block_in_R3_C2_dqdPE2(minv_block_in_R3_C2_dqdPE2) enable((*inhigh*) EN_minv_block_in_R3_C2_dqdPE2) ;
    method minv_block_in_R4_C2_dqdPE2(minv_block_in_R4_C2_dqdPE2) enable((*inhigh*) EN_minv_block_in_R4_C2_dqdPE2) ;
    method minv_block_in_R5_C2_dqdPE2(minv_block_in_R5_C2_dqdPE2) enable((*inhigh*) EN_minv_block_in_R5_C2_dqdPE2) ;
    method minv_block_in_R6_C2_dqdPE2(minv_block_in_R6_C2_dqdPE2) enable((*inhigh*) EN_minv_block_in_R6_C2_dqdPE2) ;
    method minv_block_in_R7_C2_dqdPE2(minv_block_in_R7_C2_dqdPE2) enable((*inhigh*) EN_minv_block_in_R7_C2_dqdPE2) ;
    method minv_block_in_R1_C3_dqdPE2(minv_block_in_R1_C3_dqdPE2) enable((*inhigh*) EN_minv_block_in_R1_C3_dqdPE2) ;
    method minv_block_in_R2_C3_dqdPE2(minv_block_in_R2_C3_dqdPE2) enable((*inhigh*) EN_minv_block_in_R2_C3_dqdPE2) ;
    method minv_block_in_R3_C3_dqdPE2(minv_block_in_R3_C3_dqdPE2) enable((*inhigh*) EN_minv_block_in_R3_C3_dqdPE2) ;
    method minv_block_in_R4_C3_dqdPE2(minv_block_in_R4_C3_dqdPE2) enable((*inhigh*) EN_minv_block_in_R4_C3_dqdPE2) ;
    method minv_block_in_R5_C3_dqdPE2(minv_block_in_R5_C3_dqdPE2) enable((*inhigh*) EN_minv_block_in_R5_C3_dqdPE2) ;
    method minv_block_in_R6_C3_dqdPE2(minv_block_in_R6_C3_dqdPE2) enable((*inhigh*) EN_minv_block_in_R6_C3_dqdPE2) ;
    method minv_block_in_R7_C3_dqdPE2(minv_block_in_R7_C3_dqdPE2) enable((*inhigh*) EN_minv_block_in_R7_C3_dqdPE2) ;
    method minv_block_in_R1_C4_dqdPE2(minv_block_in_R1_C4_dqdPE2) enable((*inhigh*) EN_minv_block_in_R1_C4_dqdPE2) ;
    method minv_block_in_R2_C4_dqdPE2(minv_block_in_R2_C4_dqdPE2) enable((*inhigh*) EN_minv_block_in_R2_C4_dqdPE2) ;
    method minv_block_in_R3_C4_dqdPE2(minv_block_in_R3_C4_dqdPE2) enable((*inhigh*) EN_minv_block_in_R3_C4_dqdPE2) ;
    method minv_block_in_R4_C4_dqdPE2(minv_block_in_R4_C4_dqdPE2) enable((*inhigh*) EN_minv_block_in_R4_C4_dqdPE2) ;
    method minv_block_in_R5_C4_dqdPE2(minv_block_in_R5_C4_dqdPE2) enable((*inhigh*) EN_minv_block_in_R5_C4_dqdPE2) ;
    method minv_block_in_R6_C4_dqdPE2(minv_block_in_R6_C4_dqdPE2) enable((*inhigh*) EN_minv_block_in_R6_C4_dqdPE2) ;
    method minv_block_in_R7_C4_dqdPE2(minv_block_in_R7_C4_dqdPE2) enable((*inhigh*) EN_minv_block_in_R7_C4_dqdPE2) ;
    method minv_block_in_R1_C5_dqdPE2(minv_block_in_R1_C5_dqdPE2) enable((*inhigh*) EN_minv_block_in_R1_C5_dqdPE2) ;
    method minv_block_in_R2_C5_dqdPE2(minv_block_in_R2_C5_dqdPE2) enable((*inhigh*) EN_minv_block_in_R2_C5_dqdPE2) ;
    method minv_block_in_R3_C5_dqdPE2(minv_block_in_R3_C5_dqdPE2) enable((*inhigh*) EN_minv_block_in_R3_C5_dqdPE2) ;
    method minv_block_in_R4_C5_dqdPE2(minv_block_in_R4_C5_dqdPE2) enable((*inhigh*) EN_minv_block_in_R4_C5_dqdPE2) ;
    method minv_block_in_R5_C5_dqdPE2(minv_block_in_R5_C5_dqdPE2) enable((*inhigh*) EN_minv_block_in_R5_C5_dqdPE2) ;
    method minv_block_in_R6_C5_dqdPE2(minv_block_in_R6_C5_dqdPE2) enable((*inhigh*) EN_minv_block_in_R6_C5_dqdPE2) ;
    method minv_block_in_R7_C5_dqdPE2(minv_block_in_R7_C5_dqdPE2) enable((*inhigh*) EN_minv_block_in_R7_C5_dqdPE2) ;
    method minv_block_in_R1_C6_dqdPE2(minv_block_in_R1_C6_dqdPE2) enable((*inhigh*) EN_minv_block_in_R1_C6_dqdPE2) ;
    method minv_block_in_R2_C6_dqdPE2(minv_block_in_R2_C6_dqdPE2) enable((*inhigh*) EN_minv_block_in_R2_C6_dqdPE2) ;
    method minv_block_in_R3_C6_dqdPE2(minv_block_in_R3_C6_dqdPE2) enable((*inhigh*) EN_minv_block_in_R3_C6_dqdPE2) ;
    method minv_block_in_R4_C6_dqdPE2(minv_block_in_R4_C6_dqdPE2) enable((*inhigh*) EN_minv_block_in_R4_C6_dqdPE2) ;
    method minv_block_in_R5_C6_dqdPE2(minv_block_in_R5_C6_dqdPE2) enable((*inhigh*) EN_minv_block_in_R5_C6_dqdPE2) ;
    method minv_block_in_R6_C6_dqdPE2(minv_block_in_R6_C6_dqdPE2) enable((*inhigh*) EN_minv_block_in_R6_C6_dqdPE2) ;
    method minv_block_in_R7_C6_dqdPE2(minv_block_in_R7_C6_dqdPE2) enable((*inhigh*) EN_minv_block_in_R7_C6_dqdPE2) ;
    method minv_block_in_R1_C7_dqdPE2(minv_block_in_R1_C7_dqdPE2) enable((*inhigh*) EN_minv_block_in_R1_C7_dqdPE2) ;
    method minv_block_in_R2_C7_dqdPE2(minv_block_in_R2_C7_dqdPE2) enable((*inhigh*) EN_minv_block_in_R2_C7_dqdPE2) ;
    method minv_block_in_R3_C7_dqdPE2(minv_block_in_R3_C7_dqdPE2) enable((*inhigh*) EN_minv_block_in_R3_C7_dqdPE2) ;
    method minv_block_in_R4_C7_dqdPE2(minv_block_in_R4_C7_dqdPE2) enable((*inhigh*) EN_minv_block_in_R4_C7_dqdPE2) ;
    method minv_block_in_R5_C7_dqdPE2(minv_block_in_R5_C7_dqdPE2) enable((*inhigh*) EN_minv_block_in_R5_C7_dqdPE2) ;
    method minv_block_in_R6_C7_dqdPE2(minv_block_in_R6_C7_dqdPE2) enable((*inhigh*) EN_minv_block_in_R6_C7_dqdPE2) ;
    method minv_block_in_R7_C7_dqdPE2(minv_block_in_R7_C7_dqdPE2) enable((*inhigh*) EN_minv_block_in_R7_C7_dqdPE2) ;
    method minv_block_in_R1_C1_dqdPE3(minv_block_in_R1_C1_dqdPE3) enable((*inhigh*) EN_minv_block_in_R1_C1_dqdPE3) ;
    method minv_block_in_R2_C1_dqdPE3(minv_block_in_R2_C1_dqdPE3) enable((*inhigh*) EN_minv_block_in_R2_C1_dqdPE3) ;
    method minv_block_in_R3_C1_dqdPE3(minv_block_in_R3_C1_dqdPE3) enable((*inhigh*) EN_minv_block_in_R3_C1_dqdPE3) ;
    method minv_block_in_R4_C1_dqdPE3(minv_block_in_R4_C1_dqdPE3) enable((*inhigh*) EN_minv_block_in_R4_C1_dqdPE3) ;
    method minv_block_in_R5_C1_dqdPE3(minv_block_in_R5_C1_dqdPE3) enable((*inhigh*) EN_minv_block_in_R5_C1_dqdPE3) ;
    method minv_block_in_R6_C1_dqdPE3(minv_block_in_R6_C1_dqdPE3) enable((*inhigh*) EN_minv_block_in_R6_C1_dqdPE3) ;
    method minv_block_in_R7_C1_dqdPE3(minv_block_in_R7_C1_dqdPE3) enable((*inhigh*) EN_minv_block_in_R7_C1_dqdPE3) ;
    method minv_block_in_R1_C2_dqdPE3(minv_block_in_R1_C2_dqdPE3) enable((*inhigh*) EN_minv_block_in_R1_C2_dqdPE3) ;
    method minv_block_in_R2_C2_dqdPE3(minv_block_in_R2_C2_dqdPE3) enable((*inhigh*) EN_minv_block_in_R2_C2_dqdPE3) ;
    method minv_block_in_R3_C2_dqdPE3(minv_block_in_R3_C2_dqdPE3) enable((*inhigh*) EN_minv_block_in_R3_C2_dqdPE3) ;
    method minv_block_in_R4_C2_dqdPE3(minv_block_in_R4_C2_dqdPE3) enable((*inhigh*) EN_minv_block_in_R4_C2_dqdPE3) ;
    method minv_block_in_R5_C2_dqdPE3(minv_block_in_R5_C2_dqdPE3) enable((*inhigh*) EN_minv_block_in_R5_C2_dqdPE3) ;
    method minv_block_in_R6_C2_dqdPE3(minv_block_in_R6_C2_dqdPE3) enable((*inhigh*) EN_minv_block_in_R6_C2_dqdPE3) ;
    method minv_block_in_R7_C2_dqdPE3(minv_block_in_R7_C2_dqdPE3) enable((*inhigh*) EN_minv_block_in_R7_C2_dqdPE3) ;
    method minv_block_in_R1_C3_dqdPE3(minv_block_in_R1_C3_dqdPE3) enable((*inhigh*) EN_minv_block_in_R1_C3_dqdPE3) ;
    method minv_block_in_R2_C3_dqdPE3(minv_block_in_R2_C3_dqdPE3) enable((*inhigh*) EN_minv_block_in_R2_C3_dqdPE3) ;
    method minv_block_in_R3_C3_dqdPE3(minv_block_in_R3_C3_dqdPE3) enable((*inhigh*) EN_minv_block_in_R3_C3_dqdPE3) ;
    method minv_block_in_R4_C3_dqdPE3(minv_block_in_R4_C3_dqdPE3) enable((*inhigh*) EN_minv_block_in_R4_C3_dqdPE3) ;
    method minv_block_in_R5_C3_dqdPE3(minv_block_in_R5_C3_dqdPE3) enable((*inhigh*) EN_minv_block_in_R5_C3_dqdPE3) ;
    method minv_block_in_R6_C3_dqdPE3(minv_block_in_R6_C3_dqdPE3) enable((*inhigh*) EN_minv_block_in_R6_C3_dqdPE3) ;
    method minv_block_in_R7_C3_dqdPE3(minv_block_in_R7_C3_dqdPE3) enable((*inhigh*) EN_minv_block_in_R7_C3_dqdPE3) ;
    method minv_block_in_R1_C4_dqdPE3(minv_block_in_R1_C4_dqdPE3) enable((*inhigh*) EN_minv_block_in_R1_C4_dqdPE3) ;
    method minv_block_in_R2_C4_dqdPE3(minv_block_in_R2_C4_dqdPE3) enable((*inhigh*) EN_minv_block_in_R2_C4_dqdPE3) ;
    method minv_block_in_R3_C4_dqdPE3(minv_block_in_R3_C4_dqdPE3) enable((*inhigh*) EN_minv_block_in_R3_C4_dqdPE3) ;
    method minv_block_in_R4_C4_dqdPE3(minv_block_in_R4_C4_dqdPE3) enable((*inhigh*) EN_minv_block_in_R4_C4_dqdPE3) ;
    method minv_block_in_R5_C4_dqdPE3(minv_block_in_R5_C4_dqdPE3) enable((*inhigh*) EN_minv_block_in_R5_C4_dqdPE3) ;
    method minv_block_in_R6_C4_dqdPE3(minv_block_in_R6_C4_dqdPE3) enable((*inhigh*) EN_minv_block_in_R6_C4_dqdPE3) ;
    method minv_block_in_R7_C4_dqdPE3(minv_block_in_R7_C4_dqdPE3) enable((*inhigh*) EN_minv_block_in_R7_C4_dqdPE3) ;
    method minv_block_in_R1_C5_dqdPE3(minv_block_in_R1_C5_dqdPE3) enable((*inhigh*) EN_minv_block_in_R1_C5_dqdPE3) ;
    method minv_block_in_R2_C5_dqdPE3(minv_block_in_R2_C5_dqdPE3) enable((*inhigh*) EN_minv_block_in_R2_C5_dqdPE3) ;
    method minv_block_in_R3_C5_dqdPE3(minv_block_in_R3_C5_dqdPE3) enable((*inhigh*) EN_minv_block_in_R3_C5_dqdPE3) ;
    method minv_block_in_R4_C5_dqdPE3(minv_block_in_R4_C5_dqdPE3) enable((*inhigh*) EN_minv_block_in_R4_C5_dqdPE3) ;
    method minv_block_in_R5_C5_dqdPE3(minv_block_in_R5_C5_dqdPE3) enable((*inhigh*) EN_minv_block_in_R5_C5_dqdPE3) ;
    method minv_block_in_R6_C5_dqdPE3(minv_block_in_R6_C5_dqdPE3) enable((*inhigh*) EN_minv_block_in_R6_C5_dqdPE3) ;
    method minv_block_in_R7_C5_dqdPE3(minv_block_in_R7_C5_dqdPE3) enable((*inhigh*) EN_minv_block_in_R7_C5_dqdPE3) ;
    method minv_block_in_R1_C6_dqdPE3(minv_block_in_R1_C6_dqdPE3) enable((*inhigh*) EN_minv_block_in_R1_C6_dqdPE3) ;
    method minv_block_in_R2_C6_dqdPE3(minv_block_in_R2_C6_dqdPE3) enable((*inhigh*) EN_minv_block_in_R2_C6_dqdPE3) ;
    method minv_block_in_R3_C6_dqdPE3(minv_block_in_R3_C6_dqdPE3) enable((*inhigh*) EN_minv_block_in_R3_C6_dqdPE3) ;
    method minv_block_in_R4_C6_dqdPE3(minv_block_in_R4_C6_dqdPE3) enable((*inhigh*) EN_minv_block_in_R4_C6_dqdPE3) ;
    method minv_block_in_R5_C6_dqdPE3(minv_block_in_R5_C6_dqdPE3) enable((*inhigh*) EN_minv_block_in_R5_C6_dqdPE3) ;
    method minv_block_in_R6_C6_dqdPE3(minv_block_in_R6_C6_dqdPE3) enable((*inhigh*) EN_minv_block_in_R6_C6_dqdPE3) ;
    method minv_block_in_R7_C6_dqdPE3(minv_block_in_R7_C6_dqdPE3) enable((*inhigh*) EN_minv_block_in_R7_C6_dqdPE3) ;
    method minv_block_in_R1_C7_dqdPE3(minv_block_in_R1_C7_dqdPE3) enable((*inhigh*) EN_minv_block_in_R1_C7_dqdPE3) ;
    method minv_block_in_R2_C7_dqdPE3(minv_block_in_R2_C7_dqdPE3) enable((*inhigh*) EN_minv_block_in_R2_C7_dqdPE3) ;
    method minv_block_in_R3_C7_dqdPE3(minv_block_in_R3_C7_dqdPE3) enable((*inhigh*) EN_minv_block_in_R3_C7_dqdPE3) ;
    method minv_block_in_R4_C7_dqdPE3(minv_block_in_R4_C7_dqdPE3) enable((*inhigh*) EN_minv_block_in_R4_C7_dqdPE3) ;
    method minv_block_in_R5_C7_dqdPE3(minv_block_in_R5_C7_dqdPE3) enable((*inhigh*) EN_minv_block_in_R5_C7_dqdPE3) ;
    method minv_block_in_R6_C7_dqdPE3(minv_block_in_R6_C7_dqdPE3) enable((*inhigh*) EN_minv_block_in_R6_C7_dqdPE3) ;
    method minv_block_in_R7_C7_dqdPE3(minv_block_in_R7_C7_dqdPE3) enable((*inhigh*) EN_minv_block_in_R7_C7_dqdPE3) ;
    method minv_block_in_R1_C1_dqdPE4(minv_block_in_R1_C1_dqdPE4) enable((*inhigh*) EN_minv_block_in_R1_C1_dqdPE4) ;
    method minv_block_in_R2_C1_dqdPE4(minv_block_in_R2_C1_dqdPE4) enable((*inhigh*) EN_minv_block_in_R2_C1_dqdPE4) ;
    method minv_block_in_R3_C1_dqdPE4(minv_block_in_R3_C1_dqdPE4) enable((*inhigh*) EN_minv_block_in_R3_C1_dqdPE4) ;
    method minv_block_in_R4_C1_dqdPE4(minv_block_in_R4_C1_dqdPE4) enable((*inhigh*) EN_minv_block_in_R4_C1_dqdPE4) ;
    method minv_block_in_R5_C1_dqdPE4(minv_block_in_R5_C1_dqdPE4) enable((*inhigh*) EN_minv_block_in_R5_C1_dqdPE4) ;
    method minv_block_in_R6_C1_dqdPE4(minv_block_in_R6_C1_dqdPE4) enable((*inhigh*) EN_minv_block_in_R6_C1_dqdPE4) ;
    method minv_block_in_R7_C1_dqdPE4(minv_block_in_R7_C1_dqdPE4) enable((*inhigh*) EN_minv_block_in_R7_C1_dqdPE4) ;
    method minv_block_in_R1_C2_dqdPE4(minv_block_in_R1_C2_dqdPE4) enable((*inhigh*) EN_minv_block_in_R1_C2_dqdPE4) ;
    method minv_block_in_R2_C2_dqdPE4(minv_block_in_R2_C2_dqdPE4) enable((*inhigh*) EN_minv_block_in_R2_C2_dqdPE4) ;
    method minv_block_in_R3_C2_dqdPE4(minv_block_in_R3_C2_dqdPE4) enable((*inhigh*) EN_minv_block_in_R3_C2_dqdPE4) ;
    method minv_block_in_R4_C2_dqdPE4(minv_block_in_R4_C2_dqdPE4) enable((*inhigh*) EN_minv_block_in_R4_C2_dqdPE4) ;
    method minv_block_in_R5_C2_dqdPE4(minv_block_in_R5_C2_dqdPE4) enable((*inhigh*) EN_minv_block_in_R5_C2_dqdPE4) ;
    method minv_block_in_R6_C2_dqdPE4(minv_block_in_R6_C2_dqdPE4) enable((*inhigh*) EN_minv_block_in_R6_C2_dqdPE4) ;
    method minv_block_in_R7_C2_dqdPE4(minv_block_in_R7_C2_dqdPE4) enable((*inhigh*) EN_minv_block_in_R7_C2_dqdPE4) ;
    method minv_block_in_R1_C3_dqdPE4(minv_block_in_R1_C3_dqdPE4) enable((*inhigh*) EN_minv_block_in_R1_C3_dqdPE4) ;
    method minv_block_in_R2_C3_dqdPE4(minv_block_in_R2_C3_dqdPE4) enable((*inhigh*) EN_minv_block_in_R2_C3_dqdPE4) ;
    method minv_block_in_R3_C3_dqdPE4(minv_block_in_R3_C3_dqdPE4) enable((*inhigh*) EN_minv_block_in_R3_C3_dqdPE4) ;
    method minv_block_in_R4_C3_dqdPE4(minv_block_in_R4_C3_dqdPE4) enable((*inhigh*) EN_minv_block_in_R4_C3_dqdPE4) ;
    method minv_block_in_R5_C3_dqdPE4(minv_block_in_R5_C3_dqdPE4) enable((*inhigh*) EN_minv_block_in_R5_C3_dqdPE4) ;
    method minv_block_in_R6_C3_dqdPE4(minv_block_in_R6_C3_dqdPE4) enable((*inhigh*) EN_minv_block_in_R6_C3_dqdPE4) ;
    method minv_block_in_R7_C3_dqdPE4(minv_block_in_R7_C3_dqdPE4) enable((*inhigh*) EN_minv_block_in_R7_C3_dqdPE4) ;
    method minv_block_in_R1_C4_dqdPE4(minv_block_in_R1_C4_dqdPE4) enable((*inhigh*) EN_minv_block_in_R1_C4_dqdPE4) ;
    method minv_block_in_R2_C4_dqdPE4(minv_block_in_R2_C4_dqdPE4) enable((*inhigh*) EN_minv_block_in_R2_C4_dqdPE4) ;
    method minv_block_in_R3_C4_dqdPE4(minv_block_in_R3_C4_dqdPE4) enable((*inhigh*) EN_minv_block_in_R3_C4_dqdPE4) ;
    method minv_block_in_R4_C4_dqdPE4(minv_block_in_R4_C4_dqdPE4) enable((*inhigh*) EN_minv_block_in_R4_C4_dqdPE4) ;
    method minv_block_in_R5_C4_dqdPE4(minv_block_in_R5_C4_dqdPE4) enable((*inhigh*) EN_minv_block_in_R5_C4_dqdPE4) ;
    method minv_block_in_R6_C4_dqdPE4(minv_block_in_R6_C4_dqdPE4) enable((*inhigh*) EN_minv_block_in_R6_C4_dqdPE4) ;
    method minv_block_in_R7_C4_dqdPE4(minv_block_in_R7_C4_dqdPE4) enable((*inhigh*) EN_minv_block_in_R7_C4_dqdPE4) ;
    method minv_block_in_R1_C5_dqdPE4(minv_block_in_R1_C5_dqdPE4) enable((*inhigh*) EN_minv_block_in_R1_C5_dqdPE4) ;
    method minv_block_in_R2_C5_dqdPE4(minv_block_in_R2_C5_dqdPE4) enable((*inhigh*) EN_minv_block_in_R2_C5_dqdPE4) ;
    method minv_block_in_R3_C5_dqdPE4(minv_block_in_R3_C5_dqdPE4) enable((*inhigh*) EN_minv_block_in_R3_C5_dqdPE4) ;
    method minv_block_in_R4_C5_dqdPE4(minv_block_in_R4_C5_dqdPE4) enable((*inhigh*) EN_minv_block_in_R4_C5_dqdPE4) ;
    method minv_block_in_R5_C5_dqdPE4(minv_block_in_R5_C5_dqdPE4) enable((*inhigh*) EN_minv_block_in_R5_C5_dqdPE4) ;
    method minv_block_in_R6_C5_dqdPE4(minv_block_in_R6_C5_dqdPE4) enable((*inhigh*) EN_minv_block_in_R6_C5_dqdPE4) ;
    method minv_block_in_R7_C5_dqdPE4(minv_block_in_R7_C5_dqdPE4) enable((*inhigh*) EN_minv_block_in_R7_C5_dqdPE4) ;
    method minv_block_in_R1_C6_dqdPE4(minv_block_in_R1_C6_dqdPE4) enable((*inhigh*) EN_minv_block_in_R1_C6_dqdPE4) ;
    method minv_block_in_R2_C6_dqdPE4(minv_block_in_R2_C6_dqdPE4) enable((*inhigh*) EN_minv_block_in_R2_C6_dqdPE4) ;
    method minv_block_in_R3_C6_dqdPE4(minv_block_in_R3_C6_dqdPE4) enable((*inhigh*) EN_minv_block_in_R3_C6_dqdPE4) ;
    method minv_block_in_R4_C6_dqdPE4(minv_block_in_R4_C6_dqdPE4) enable((*inhigh*) EN_minv_block_in_R4_C6_dqdPE4) ;
    method minv_block_in_R5_C6_dqdPE4(minv_block_in_R5_C6_dqdPE4) enable((*inhigh*) EN_minv_block_in_R5_C6_dqdPE4) ;
    method minv_block_in_R6_C6_dqdPE4(minv_block_in_R6_C6_dqdPE4) enable((*inhigh*) EN_minv_block_in_R6_C6_dqdPE4) ;
    method minv_block_in_R7_C6_dqdPE4(minv_block_in_R7_C6_dqdPE4) enable((*inhigh*) EN_minv_block_in_R7_C6_dqdPE4) ;
    method minv_block_in_R1_C7_dqdPE4(minv_block_in_R1_C7_dqdPE4) enable((*inhigh*) EN_minv_block_in_R1_C7_dqdPE4) ;
    method minv_block_in_R2_C7_dqdPE4(minv_block_in_R2_C7_dqdPE4) enable((*inhigh*) EN_minv_block_in_R2_C7_dqdPE4) ;
    method minv_block_in_R3_C7_dqdPE4(minv_block_in_R3_C7_dqdPE4) enable((*inhigh*) EN_minv_block_in_R3_C7_dqdPE4) ;
    method minv_block_in_R4_C7_dqdPE4(minv_block_in_R4_C7_dqdPE4) enable((*inhigh*) EN_minv_block_in_R4_C7_dqdPE4) ;
    method minv_block_in_R5_C7_dqdPE4(minv_block_in_R5_C7_dqdPE4) enable((*inhigh*) EN_minv_block_in_R5_C7_dqdPE4) ;
    method minv_block_in_R6_C7_dqdPE4(minv_block_in_R6_C7_dqdPE4) enable((*inhigh*) EN_minv_block_in_R6_C7_dqdPE4) ;
    method minv_block_in_R7_C7_dqdPE4(minv_block_in_R7_C7_dqdPE4) enable((*inhigh*) EN_minv_block_in_R7_C7_dqdPE4) ;
    method minv_block_in_R1_C1_dqdPE5(minv_block_in_R1_C1_dqdPE5) enable((*inhigh*) EN_minv_block_in_R1_C1_dqdPE5) ;
    method minv_block_in_R2_C1_dqdPE5(minv_block_in_R2_C1_dqdPE5) enable((*inhigh*) EN_minv_block_in_R2_C1_dqdPE5) ;
    method minv_block_in_R3_C1_dqdPE5(minv_block_in_R3_C1_dqdPE5) enable((*inhigh*) EN_minv_block_in_R3_C1_dqdPE5) ;
    method minv_block_in_R4_C1_dqdPE5(minv_block_in_R4_C1_dqdPE5) enable((*inhigh*) EN_minv_block_in_R4_C1_dqdPE5) ;
    method minv_block_in_R5_C1_dqdPE5(minv_block_in_R5_C1_dqdPE5) enable((*inhigh*) EN_minv_block_in_R5_C1_dqdPE5) ;
    method minv_block_in_R6_C1_dqdPE5(minv_block_in_R6_C1_dqdPE5) enable((*inhigh*) EN_minv_block_in_R6_C1_dqdPE5) ;
    method minv_block_in_R7_C1_dqdPE5(minv_block_in_R7_C1_dqdPE5) enable((*inhigh*) EN_minv_block_in_R7_C1_dqdPE5) ;
    method minv_block_in_R1_C2_dqdPE5(minv_block_in_R1_C2_dqdPE5) enable((*inhigh*) EN_minv_block_in_R1_C2_dqdPE5) ;
    method minv_block_in_R2_C2_dqdPE5(minv_block_in_R2_C2_dqdPE5) enable((*inhigh*) EN_minv_block_in_R2_C2_dqdPE5) ;
    method minv_block_in_R3_C2_dqdPE5(minv_block_in_R3_C2_dqdPE5) enable((*inhigh*) EN_minv_block_in_R3_C2_dqdPE5) ;
    method minv_block_in_R4_C2_dqdPE5(minv_block_in_R4_C2_dqdPE5) enable((*inhigh*) EN_minv_block_in_R4_C2_dqdPE5) ;
    method minv_block_in_R5_C2_dqdPE5(minv_block_in_R5_C2_dqdPE5) enable((*inhigh*) EN_minv_block_in_R5_C2_dqdPE5) ;
    method minv_block_in_R6_C2_dqdPE5(minv_block_in_R6_C2_dqdPE5) enable((*inhigh*) EN_minv_block_in_R6_C2_dqdPE5) ;
    method minv_block_in_R7_C2_dqdPE5(minv_block_in_R7_C2_dqdPE5) enable((*inhigh*) EN_minv_block_in_R7_C2_dqdPE5) ;
    method minv_block_in_R1_C3_dqdPE5(minv_block_in_R1_C3_dqdPE5) enable((*inhigh*) EN_minv_block_in_R1_C3_dqdPE5) ;
    method minv_block_in_R2_C3_dqdPE5(minv_block_in_R2_C3_dqdPE5) enable((*inhigh*) EN_minv_block_in_R2_C3_dqdPE5) ;
    method minv_block_in_R3_C3_dqdPE5(minv_block_in_R3_C3_dqdPE5) enable((*inhigh*) EN_minv_block_in_R3_C3_dqdPE5) ;
    method minv_block_in_R4_C3_dqdPE5(minv_block_in_R4_C3_dqdPE5) enable((*inhigh*) EN_minv_block_in_R4_C3_dqdPE5) ;
    method minv_block_in_R5_C3_dqdPE5(minv_block_in_R5_C3_dqdPE5) enable((*inhigh*) EN_minv_block_in_R5_C3_dqdPE5) ;
    method minv_block_in_R6_C3_dqdPE5(minv_block_in_R6_C3_dqdPE5) enable((*inhigh*) EN_minv_block_in_R6_C3_dqdPE5) ;
    method minv_block_in_R7_C3_dqdPE5(minv_block_in_R7_C3_dqdPE5) enable((*inhigh*) EN_minv_block_in_R7_C3_dqdPE5) ;
    method minv_block_in_R1_C4_dqdPE5(minv_block_in_R1_C4_dqdPE5) enable((*inhigh*) EN_minv_block_in_R1_C4_dqdPE5) ;
    method minv_block_in_R2_C4_dqdPE5(minv_block_in_R2_C4_dqdPE5) enable((*inhigh*) EN_minv_block_in_R2_C4_dqdPE5) ;
    method minv_block_in_R3_C4_dqdPE5(minv_block_in_R3_C4_dqdPE5) enable((*inhigh*) EN_minv_block_in_R3_C4_dqdPE5) ;
    method minv_block_in_R4_C4_dqdPE5(minv_block_in_R4_C4_dqdPE5) enable((*inhigh*) EN_minv_block_in_R4_C4_dqdPE5) ;
    method minv_block_in_R5_C4_dqdPE5(minv_block_in_R5_C4_dqdPE5) enable((*inhigh*) EN_minv_block_in_R5_C4_dqdPE5) ;
    method minv_block_in_R6_C4_dqdPE5(minv_block_in_R6_C4_dqdPE5) enable((*inhigh*) EN_minv_block_in_R6_C4_dqdPE5) ;
    method minv_block_in_R7_C4_dqdPE5(minv_block_in_R7_C4_dqdPE5) enable((*inhigh*) EN_minv_block_in_R7_C4_dqdPE5) ;
    method minv_block_in_R1_C5_dqdPE5(minv_block_in_R1_C5_dqdPE5) enable((*inhigh*) EN_minv_block_in_R1_C5_dqdPE5) ;
    method minv_block_in_R2_C5_dqdPE5(minv_block_in_R2_C5_dqdPE5) enable((*inhigh*) EN_minv_block_in_R2_C5_dqdPE5) ;
    method minv_block_in_R3_C5_dqdPE5(minv_block_in_R3_C5_dqdPE5) enable((*inhigh*) EN_minv_block_in_R3_C5_dqdPE5) ;
    method minv_block_in_R4_C5_dqdPE5(minv_block_in_R4_C5_dqdPE5) enable((*inhigh*) EN_minv_block_in_R4_C5_dqdPE5) ;
    method minv_block_in_R5_C5_dqdPE5(minv_block_in_R5_C5_dqdPE5) enable((*inhigh*) EN_minv_block_in_R5_C5_dqdPE5) ;
    method minv_block_in_R6_C5_dqdPE5(minv_block_in_R6_C5_dqdPE5) enable((*inhigh*) EN_minv_block_in_R6_C5_dqdPE5) ;
    method minv_block_in_R7_C5_dqdPE5(minv_block_in_R7_C5_dqdPE5) enable((*inhigh*) EN_minv_block_in_R7_C5_dqdPE5) ;
    method minv_block_in_R1_C6_dqdPE5(minv_block_in_R1_C6_dqdPE5) enable((*inhigh*) EN_minv_block_in_R1_C6_dqdPE5) ;
    method minv_block_in_R2_C6_dqdPE5(minv_block_in_R2_C6_dqdPE5) enable((*inhigh*) EN_minv_block_in_R2_C6_dqdPE5) ;
    method minv_block_in_R3_C6_dqdPE5(minv_block_in_R3_C6_dqdPE5) enable((*inhigh*) EN_minv_block_in_R3_C6_dqdPE5) ;
    method minv_block_in_R4_C6_dqdPE5(minv_block_in_R4_C6_dqdPE5) enable((*inhigh*) EN_minv_block_in_R4_C6_dqdPE5) ;
    method minv_block_in_R5_C6_dqdPE5(minv_block_in_R5_C6_dqdPE5) enable((*inhigh*) EN_minv_block_in_R5_C6_dqdPE5) ;
    method minv_block_in_R6_C6_dqdPE5(minv_block_in_R6_C6_dqdPE5) enable((*inhigh*) EN_minv_block_in_R6_C6_dqdPE5) ;
    method minv_block_in_R7_C6_dqdPE5(minv_block_in_R7_C6_dqdPE5) enable((*inhigh*) EN_minv_block_in_R7_C6_dqdPE5) ;
    method minv_block_in_R1_C7_dqdPE5(minv_block_in_R1_C7_dqdPE5) enable((*inhigh*) EN_minv_block_in_R1_C7_dqdPE5) ;
    method minv_block_in_R2_C7_dqdPE5(minv_block_in_R2_C7_dqdPE5) enable((*inhigh*) EN_minv_block_in_R2_C7_dqdPE5) ;
    method minv_block_in_R3_C7_dqdPE5(minv_block_in_R3_C7_dqdPE5) enable((*inhigh*) EN_minv_block_in_R3_C7_dqdPE5) ;
    method minv_block_in_R4_C7_dqdPE5(minv_block_in_R4_C7_dqdPE5) enable((*inhigh*) EN_minv_block_in_R4_C7_dqdPE5) ;
    method minv_block_in_R5_C7_dqdPE5(minv_block_in_R5_C7_dqdPE5) enable((*inhigh*) EN_minv_block_in_R5_C7_dqdPE5) ;
    method minv_block_in_R6_C7_dqdPE5(minv_block_in_R6_C7_dqdPE5) enable((*inhigh*) EN_minv_block_in_R6_C7_dqdPE5) ;
    method minv_block_in_R7_C7_dqdPE5(minv_block_in_R7_C7_dqdPE5) enable((*inhigh*) EN_minv_block_in_R7_C7_dqdPE5) ;
    method minv_block_in_R1_C1_dqdPE6(minv_block_in_R1_C1_dqdPE6) enable((*inhigh*) EN_minv_block_in_R1_C1_dqdPE6) ;
    method minv_block_in_R2_C1_dqdPE6(minv_block_in_R2_C1_dqdPE6) enable((*inhigh*) EN_minv_block_in_R2_C1_dqdPE6) ;
    method minv_block_in_R3_C1_dqdPE6(minv_block_in_R3_C1_dqdPE6) enable((*inhigh*) EN_minv_block_in_R3_C1_dqdPE6) ;
    method minv_block_in_R4_C1_dqdPE6(minv_block_in_R4_C1_dqdPE6) enable((*inhigh*) EN_minv_block_in_R4_C1_dqdPE6) ;
    method minv_block_in_R5_C1_dqdPE6(minv_block_in_R5_C1_dqdPE6) enable((*inhigh*) EN_minv_block_in_R5_C1_dqdPE6) ;
    method minv_block_in_R6_C1_dqdPE6(minv_block_in_R6_C1_dqdPE6) enable((*inhigh*) EN_minv_block_in_R6_C1_dqdPE6) ;
    method minv_block_in_R7_C1_dqdPE6(minv_block_in_R7_C1_dqdPE6) enable((*inhigh*) EN_minv_block_in_R7_C1_dqdPE6) ;
    method minv_block_in_R1_C2_dqdPE6(minv_block_in_R1_C2_dqdPE6) enable((*inhigh*) EN_minv_block_in_R1_C2_dqdPE6) ;
    method minv_block_in_R2_C2_dqdPE6(minv_block_in_R2_C2_dqdPE6) enable((*inhigh*) EN_minv_block_in_R2_C2_dqdPE6) ;
    method minv_block_in_R3_C2_dqdPE6(minv_block_in_R3_C2_dqdPE6) enable((*inhigh*) EN_minv_block_in_R3_C2_dqdPE6) ;
    method minv_block_in_R4_C2_dqdPE6(minv_block_in_R4_C2_dqdPE6) enable((*inhigh*) EN_minv_block_in_R4_C2_dqdPE6) ;
    method minv_block_in_R5_C2_dqdPE6(minv_block_in_R5_C2_dqdPE6) enable((*inhigh*) EN_minv_block_in_R5_C2_dqdPE6) ;
    method minv_block_in_R6_C2_dqdPE6(minv_block_in_R6_C2_dqdPE6) enable((*inhigh*) EN_minv_block_in_R6_C2_dqdPE6) ;
    method minv_block_in_R7_C2_dqdPE6(minv_block_in_R7_C2_dqdPE6) enable((*inhigh*) EN_minv_block_in_R7_C2_dqdPE6) ;
    method minv_block_in_R1_C3_dqdPE6(minv_block_in_R1_C3_dqdPE6) enable((*inhigh*) EN_minv_block_in_R1_C3_dqdPE6) ;
    method minv_block_in_R2_C3_dqdPE6(minv_block_in_R2_C3_dqdPE6) enable((*inhigh*) EN_minv_block_in_R2_C3_dqdPE6) ;
    method minv_block_in_R3_C3_dqdPE6(minv_block_in_R3_C3_dqdPE6) enable((*inhigh*) EN_minv_block_in_R3_C3_dqdPE6) ;
    method minv_block_in_R4_C3_dqdPE6(minv_block_in_R4_C3_dqdPE6) enable((*inhigh*) EN_minv_block_in_R4_C3_dqdPE6) ;
    method minv_block_in_R5_C3_dqdPE6(minv_block_in_R5_C3_dqdPE6) enable((*inhigh*) EN_minv_block_in_R5_C3_dqdPE6) ;
    method minv_block_in_R6_C3_dqdPE6(minv_block_in_R6_C3_dqdPE6) enable((*inhigh*) EN_minv_block_in_R6_C3_dqdPE6) ;
    method minv_block_in_R7_C3_dqdPE6(minv_block_in_R7_C3_dqdPE6) enable((*inhigh*) EN_minv_block_in_R7_C3_dqdPE6) ;
    method minv_block_in_R1_C4_dqdPE6(minv_block_in_R1_C4_dqdPE6) enable((*inhigh*) EN_minv_block_in_R1_C4_dqdPE6) ;
    method minv_block_in_R2_C4_dqdPE6(minv_block_in_R2_C4_dqdPE6) enable((*inhigh*) EN_minv_block_in_R2_C4_dqdPE6) ;
    method minv_block_in_R3_C4_dqdPE6(minv_block_in_R3_C4_dqdPE6) enable((*inhigh*) EN_minv_block_in_R3_C4_dqdPE6) ;
    method minv_block_in_R4_C4_dqdPE6(minv_block_in_R4_C4_dqdPE6) enable((*inhigh*) EN_minv_block_in_R4_C4_dqdPE6) ;
    method minv_block_in_R5_C4_dqdPE6(minv_block_in_R5_C4_dqdPE6) enable((*inhigh*) EN_minv_block_in_R5_C4_dqdPE6) ;
    method minv_block_in_R6_C4_dqdPE6(minv_block_in_R6_C4_dqdPE6) enable((*inhigh*) EN_minv_block_in_R6_C4_dqdPE6) ;
    method minv_block_in_R7_C4_dqdPE6(minv_block_in_R7_C4_dqdPE6) enable((*inhigh*) EN_minv_block_in_R7_C4_dqdPE6) ;
    method minv_block_in_R1_C5_dqdPE6(minv_block_in_R1_C5_dqdPE6) enable((*inhigh*) EN_minv_block_in_R1_C5_dqdPE6) ;
    method minv_block_in_R2_C5_dqdPE6(minv_block_in_R2_C5_dqdPE6) enable((*inhigh*) EN_minv_block_in_R2_C5_dqdPE6) ;
    method minv_block_in_R3_C5_dqdPE6(minv_block_in_R3_C5_dqdPE6) enable((*inhigh*) EN_minv_block_in_R3_C5_dqdPE6) ;
    method minv_block_in_R4_C5_dqdPE6(minv_block_in_R4_C5_dqdPE6) enable((*inhigh*) EN_minv_block_in_R4_C5_dqdPE6) ;
    method minv_block_in_R5_C5_dqdPE6(minv_block_in_R5_C5_dqdPE6) enable((*inhigh*) EN_minv_block_in_R5_C5_dqdPE6) ;
    method minv_block_in_R6_C5_dqdPE6(minv_block_in_R6_C5_dqdPE6) enable((*inhigh*) EN_minv_block_in_R6_C5_dqdPE6) ;
    method minv_block_in_R7_C5_dqdPE6(minv_block_in_R7_C5_dqdPE6) enable((*inhigh*) EN_minv_block_in_R7_C5_dqdPE6) ;
    method minv_block_in_R1_C6_dqdPE6(minv_block_in_R1_C6_dqdPE6) enable((*inhigh*) EN_minv_block_in_R1_C6_dqdPE6) ;
    method minv_block_in_R2_C6_dqdPE6(minv_block_in_R2_C6_dqdPE6) enable((*inhigh*) EN_minv_block_in_R2_C6_dqdPE6) ;
    method minv_block_in_R3_C6_dqdPE6(minv_block_in_R3_C6_dqdPE6) enable((*inhigh*) EN_minv_block_in_R3_C6_dqdPE6) ;
    method minv_block_in_R4_C6_dqdPE6(minv_block_in_R4_C6_dqdPE6) enable((*inhigh*) EN_minv_block_in_R4_C6_dqdPE6) ;
    method minv_block_in_R5_C6_dqdPE6(minv_block_in_R5_C6_dqdPE6) enable((*inhigh*) EN_minv_block_in_R5_C6_dqdPE6) ;
    method minv_block_in_R6_C6_dqdPE6(minv_block_in_R6_C6_dqdPE6) enable((*inhigh*) EN_minv_block_in_R6_C6_dqdPE6) ;
    method minv_block_in_R7_C6_dqdPE6(minv_block_in_R7_C6_dqdPE6) enable((*inhigh*) EN_minv_block_in_R7_C6_dqdPE6) ;
    method minv_block_in_R1_C7_dqdPE6(minv_block_in_R1_C7_dqdPE6) enable((*inhigh*) EN_minv_block_in_R1_C7_dqdPE6) ;
    method minv_block_in_R2_C7_dqdPE6(minv_block_in_R2_C7_dqdPE6) enable((*inhigh*) EN_minv_block_in_R2_C7_dqdPE6) ;
    method minv_block_in_R3_C7_dqdPE6(minv_block_in_R3_C7_dqdPE6) enable((*inhigh*) EN_minv_block_in_R3_C7_dqdPE6) ;
    method minv_block_in_R4_C7_dqdPE6(minv_block_in_R4_C7_dqdPE6) enable((*inhigh*) EN_minv_block_in_R4_C7_dqdPE6) ;
    method minv_block_in_R5_C7_dqdPE6(minv_block_in_R5_C7_dqdPE6) enable((*inhigh*) EN_minv_block_in_R5_C7_dqdPE6) ;
    method minv_block_in_R6_C7_dqdPE6(minv_block_in_R6_C7_dqdPE6) enable((*inhigh*) EN_minv_block_in_R6_C7_dqdPE6) ;
    method minv_block_in_R7_C7_dqdPE6(minv_block_in_R7_C7_dqdPE6) enable((*inhigh*) EN_minv_block_in_R7_C7_dqdPE6) ;
    method minv_block_in_R1_C1_dqdPE7(minv_block_in_R1_C1_dqdPE7) enable((*inhigh*) EN_minv_block_in_R1_C1_dqdPE7) ;
    method minv_block_in_R2_C1_dqdPE7(minv_block_in_R2_C1_dqdPE7) enable((*inhigh*) EN_minv_block_in_R2_C1_dqdPE7) ;
    method minv_block_in_R3_C1_dqdPE7(minv_block_in_R3_C1_dqdPE7) enable((*inhigh*) EN_minv_block_in_R3_C1_dqdPE7) ;
    method minv_block_in_R4_C1_dqdPE7(minv_block_in_R4_C1_dqdPE7) enable((*inhigh*) EN_minv_block_in_R4_C1_dqdPE7) ;
    method minv_block_in_R5_C1_dqdPE7(minv_block_in_R5_C1_dqdPE7) enable((*inhigh*) EN_minv_block_in_R5_C1_dqdPE7) ;
    method minv_block_in_R6_C1_dqdPE7(minv_block_in_R6_C1_dqdPE7) enable((*inhigh*) EN_minv_block_in_R6_C1_dqdPE7) ;
    method minv_block_in_R7_C1_dqdPE7(minv_block_in_R7_C1_dqdPE7) enable((*inhigh*) EN_minv_block_in_R7_C1_dqdPE7) ;
    method minv_block_in_R1_C2_dqdPE7(minv_block_in_R1_C2_dqdPE7) enable((*inhigh*) EN_minv_block_in_R1_C2_dqdPE7) ;
    method minv_block_in_R2_C2_dqdPE7(minv_block_in_R2_C2_dqdPE7) enable((*inhigh*) EN_minv_block_in_R2_C2_dqdPE7) ;
    method minv_block_in_R3_C2_dqdPE7(minv_block_in_R3_C2_dqdPE7) enable((*inhigh*) EN_minv_block_in_R3_C2_dqdPE7) ;
    method minv_block_in_R4_C2_dqdPE7(minv_block_in_R4_C2_dqdPE7) enable((*inhigh*) EN_minv_block_in_R4_C2_dqdPE7) ;
    method minv_block_in_R5_C2_dqdPE7(minv_block_in_R5_C2_dqdPE7) enable((*inhigh*) EN_minv_block_in_R5_C2_dqdPE7) ;
    method minv_block_in_R6_C2_dqdPE7(minv_block_in_R6_C2_dqdPE7) enable((*inhigh*) EN_minv_block_in_R6_C2_dqdPE7) ;
    method minv_block_in_R7_C2_dqdPE7(minv_block_in_R7_C2_dqdPE7) enable((*inhigh*) EN_minv_block_in_R7_C2_dqdPE7) ;
    method minv_block_in_R1_C3_dqdPE7(minv_block_in_R1_C3_dqdPE7) enable((*inhigh*) EN_minv_block_in_R1_C3_dqdPE7) ;
    method minv_block_in_R2_C3_dqdPE7(minv_block_in_R2_C3_dqdPE7) enable((*inhigh*) EN_minv_block_in_R2_C3_dqdPE7) ;
    method minv_block_in_R3_C3_dqdPE7(minv_block_in_R3_C3_dqdPE7) enable((*inhigh*) EN_minv_block_in_R3_C3_dqdPE7) ;
    method minv_block_in_R4_C3_dqdPE7(minv_block_in_R4_C3_dqdPE7) enable((*inhigh*) EN_minv_block_in_R4_C3_dqdPE7) ;
    method minv_block_in_R5_C3_dqdPE7(minv_block_in_R5_C3_dqdPE7) enable((*inhigh*) EN_minv_block_in_R5_C3_dqdPE7) ;
    method minv_block_in_R6_C3_dqdPE7(minv_block_in_R6_C3_dqdPE7) enable((*inhigh*) EN_minv_block_in_R6_C3_dqdPE7) ;
    method minv_block_in_R7_C3_dqdPE7(minv_block_in_R7_C3_dqdPE7) enable((*inhigh*) EN_minv_block_in_R7_C3_dqdPE7) ;
    method minv_block_in_R1_C4_dqdPE7(minv_block_in_R1_C4_dqdPE7) enable((*inhigh*) EN_minv_block_in_R1_C4_dqdPE7) ;
    method minv_block_in_R2_C4_dqdPE7(minv_block_in_R2_C4_dqdPE7) enable((*inhigh*) EN_minv_block_in_R2_C4_dqdPE7) ;
    method minv_block_in_R3_C4_dqdPE7(minv_block_in_R3_C4_dqdPE7) enable((*inhigh*) EN_minv_block_in_R3_C4_dqdPE7) ;
    method minv_block_in_R4_C4_dqdPE7(minv_block_in_R4_C4_dqdPE7) enable((*inhigh*) EN_minv_block_in_R4_C4_dqdPE7) ;
    method minv_block_in_R5_C4_dqdPE7(minv_block_in_R5_C4_dqdPE7) enable((*inhigh*) EN_minv_block_in_R5_C4_dqdPE7) ;
    method minv_block_in_R6_C4_dqdPE7(minv_block_in_R6_C4_dqdPE7) enable((*inhigh*) EN_minv_block_in_R6_C4_dqdPE7) ;
    method minv_block_in_R7_C4_dqdPE7(minv_block_in_R7_C4_dqdPE7) enable((*inhigh*) EN_minv_block_in_R7_C4_dqdPE7) ;
    method minv_block_in_R1_C5_dqdPE7(minv_block_in_R1_C5_dqdPE7) enable((*inhigh*) EN_minv_block_in_R1_C5_dqdPE7) ;
    method minv_block_in_R2_C5_dqdPE7(minv_block_in_R2_C5_dqdPE7) enable((*inhigh*) EN_minv_block_in_R2_C5_dqdPE7) ;
    method minv_block_in_R3_C5_dqdPE7(minv_block_in_R3_C5_dqdPE7) enable((*inhigh*) EN_minv_block_in_R3_C5_dqdPE7) ;
    method minv_block_in_R4_C5_dqdPE7(minv_block_in_R4_C5_dqdPE7) enable((*inhigh*) EN_minv_block_in_R4_C5_dqdPE7) ;
    method minv_block_in_R5_C5_dqdPE7(minv_block_in_R5_C5_dqdPE7) enable((*inhigh*) EN_minv_block_in_R5_C5_dqdPE7) ;
    method minv_block_in_R6_C5_dqdPE7(minv_block_in_R6_C5_dqdPE7) enable((*inhigh*) EN_minv_block_in_R6_C5_dqdPE7) ;
    method minv_block_in_R7_C5_dqdPE7(minv_block_in_R7_C5_dqdPE7) enable((*inhigh*) EN_minv_block_in_R7_C5_dqdPE7) ;
    method minv_block_in_R1_C6_dqdPE7(minv_block_in_R1_C6_dqdPE7) enable((*inhigh*) EN_minv_block_in_R1_C6_dqdPE7) ;
    method minv_block_in_R2_C6_dqdPE7(minv_block_in_R2_C6_dqdPE7) enable((*inhigh*) EN_minv_block_in_R2_C6_dqdPE7) ;
    method minv_block_in_R3_C6_dqdPE7(minv_block_in_R3_C6_dqdPE7) enable((*inhigh*) EN_minv_block_in_R3_C6_dqdPE7) ;
    method minv_block_in_R4_C6_dqdPE7(minv_block_in_R4_C6_dqdPE7) enable((*inhigh*) EN_minv_block_in_R4_C6_dqdPE7) ;
    method minv_block_in_R5_C6_dqdPE7(minv_block_in_R5_C6_dqdPE7) enable((*inhigh*) EN_minv_block_in_R5_C6_dqdPE7) ;
    method minv_block_in_R6_C6_dqdPE7(minv_block_in_R6_C6_dqdPE7) enable((*inhigh*) EN_minv_block_in_R6_C6_dqdPE7) ;
    method minv_block_in_R7_C6_dqdPE7(minv_block_in_R7_C6_dqdPE7) enable((*inhigh*) EN_minv_block_in_R7_C6_dqdPE7) ;
    method minv_block_in_R1_C7_dqdPE7(minv_block_in_R1_C7_dqdPE7) enable((*inhigh*) EN_minv_block_in_R1_C7_dqdPE7) ;
    method minv_block_in_R2_C7_dqdPE7(minv_block_in_R2_C7_dqdPE7) enable((*inhigh*) EN_minv_block_in_R2_C7_dqdPE7) ;
    method minv_block_in_R3_C7_dqdPE7(minv_block_in_R3_C7_dqdPE7) enable((*inhigh*) EN_minv_block_in_R3_C7_dqdPE7) ;
    method minv_block_in_R4_C7_dqdPE7(minv_block_in_R4_C7_dqdPE7) enable((*inhigh*) EN_minv_block_in_R4_C7_dqdPE7) ;
    method minv_block_in_R5_C7_dqdPE7(minv_block_in_R5_C7_dqdPE7) enable((*inhigh*) EN_minv_block_in_R5_C7_dqdPE7) ;
    method minv_block_in_R6_C7_dqdPE7(minv_block_in_R6_C7_dqdPE7) enable((*inhigh*) EN_minv_block_in_R6_C7_dqdPE7) ;
    method minv_block_in_R7_C7_dqdPE7(minv_block_in_R7_C7_dqdPE7) enable((*inhigh*) EN_minv_block_in_R7_C7_dqdPE7) ;
    method dtau_vec_in_R1_dqdPE1(dtau_vec_in_R1_dqdPE1) enable((*inhigh*) EN_dtau_vec_in_R1_dqdPE1) ;
    method dtau_vec_in_R2_dqdPE1(dtau_vec_in_R2_dqdPE1) enable((*inhigh*) EN_dtau_vec_in_R2_dqdPE1) ;
    method dtau_vec_in_R3_dqdPE1(dtau_vec_in_R3_dqdPE1) enable((*inhigh*) EN_dtau_vec_in_R3_dqdPE1) ;
    method dtau_vec_in_R4_dqdPE1(dtau_vec_in_R4_dqdPE1) enable((*inhigh*) EN_dtau_vec_in_R4_dqdPE1) ;
    method dtau_vec_in_R5_dqdPE1(dtau_vec_in_R5_dqdPE1) enable((*inhigh*) EN_dtau_vec_in_R5_dqdPE1) ;
    method dtau_vec_in_R6_dqdPE1(dtau_vec_in_R6_dqdPE1) enable((*inhigh*) EN_dtau_vec_in_R6_dqdPE1) ;
    method dtau_vec_in_R7_dqdPE1(dtau_vec_in_R7_dqdPE1) enable((*inhigh*) EN_dtau_vec_in_R7_dqdPE1) ;
    method dtau_vec_in_R1_dqdPE2(dtau_vec_in_R1_dqdPE2) enable((*inhigh*) EN_dtau_vec_in_R1_dqdPE2) ;
    method dtau_vec_in_R2_dqdPE2(dtau_vec_in_R2_dqdPE2) enable((*inhigh*) EN_dtau_vec_in_R2_dqdPE2) ;
    method dtau_vec_in_R3_dqdPE2(dtau_vec_in_R3_dqdPE2) enable((*inhigh*) EN_dtau_vec_in_R3_dqdPE2) ;
    method dtau_vec_in_R4_dqdPE2(dtau_vec_in_R4_dqdPE2) enable((*inhigh*) EN_dtau_vec_in_R4_dqdPE2) ;
    method dtau_vec_in_R5_dqdPE2(dtau_vec_in_R5_dqdPE2) enable((*inhigh*) EN_dtau_vec_in_R5_dqdPE2) ;
    method dtau_vec_in_R6_dqdPE2(dtau_vec_in_R6_dqdPE2) enable((*inhigh*) EN_dtau_vec_in_R6_dqdPE2) ;
    method dtau_vec_in_R7_dqdPE2(dtau_vec_in_R7_dqdPE2) enable((*inhigh*) EN_dtau_vec_in_R7_dqdPE2) ;
    method dtau_vec_in_R1_dqdPE3(dtau_vec_in_R1_dqdPE3) enable((*inhigh*) EN_dtau_vec_in_R1_dqdPE3) ;
    method dtau_vec_in_R2_dqdPE3(dtau_vec_in_R2_dqdPE3) enable((*inhigh*) EN_dtau_vec_in_R2_dqdPE3) ;
    method dtau_vec_in_R3_dqdPE3(dtau_vec_in_R3_dqdPE3) enable((*inhigh*) EN_dtau_vec_in_R3_dqdPE3) ;
    method dtau_vec_in_R4_dqdPE3(dtau_vec_in_R4_dqdPE3) enable((*inhigh*) EN_dtau_vec_in_R4_dqdPE3) ;
    method dtau_vec_in_R5_dqdPE3(dtau_vec_in_R5_dqdPE3) enable((*inhigh*) EN_dtau_vec_in_R5_dqdPE3) ;
    method dtau_vec_in_R6_dqdPE3(dtau_vec_in_R6_dqdPE3) enable((*inhigh*) EN_dtau_vec_in_R6_dqdPE3) ;
    method dtau_vec_in_R7_dqdPE3(dtau_vec_in_R7_dqdPE3) enable((*inhigh*) EN_dtau_vec_in_R7_dqdPE3) ;
    method dtau_vec_in_R1_dqdPE4(dtau_vec_in_R1_dqdPE4) enable((*inhigh*) EN_dtau_vec_in_R1_dqdPE4) ;
    method dtau_vec_in_R2_dqdPE4(dtau_vec_in_R2_dqdPE4) enable((*inhigh*) EN_dtau_vec_in_R2_dqdPE4) ;
    method dtau_vec_in_R3_dqdPE4(dtau_vec_in_R3_dqdPE4) enable((*inhigh*) EN_dtau_vec_in_R3_dqdPE4) ;
    method dtau_vec_in_R4_dqdPE4(dtau_vec_in_R4_dqdPE4) enable((*inhigh*) EN_dtau_vec_in_R4_dqdPE4) ;
    method dtau_vec_in_R5_dqdPE4(dtau_vec_in_R5_dqdPE4) enable((*inhigh*) EN_dtau_vec_in_R5_dqdPE4) ;
    method dtau_vec_in_R6_dqdPE4(dtau_vec_in_R6_dqdPE4) enable((*inhigh*) EN_dtau_vec_in_R6_dqdPE4) ;
    method dtau_vec_in_R7_dqdPE4(dtau_vec_in_R7_dqdPE4) enable((*inhigh*) EN_dtau_vec_in_R7_dqdPE4) ;
    method dtau_vec_in_R1_dqdPE5(dtau_vec_in_R1_dqdPE5) enable((*inhigh*) EN_dtau_vec_in_R1_dqdPE5) ;
    method dtau_vec_in_R2_dqdPE5(dtau_vec_in_R2_dqdPE5) enable((*inhigh*) EN_dtau_vec_in_R2_dqdPE5) ;
    method dtau_vec_in_R3_dqdPE5(dtau_vec_in_R3_dqdPE5) enable((*inhigh*) EN_dtau_vec_in_R3_dqdPE5) ;
    method dtau_vec_in_R4_dqdPE5(dtau_vec_in_R4_dqdPE5) enable((*inhigh*) EN_dtau_vec_in_R4_dqdPE5) ;
    method dtau_vec_in_R5_dqdPE5(dtau_vec_in_R5_dqdPE5) enable((*inhigh*) EN_dtau_vec_in_R5_dqdPE5) ;
    method dtau_vec_in_R6_dqdPE5(dtau_vec_in_R6_dqdPE5) enable((*inhigh*) EN_dtau_vec_in_R6_dqdPE5) ;
    method dtau_vec_in_R7_dqdPE5(dtau_vec_in_R7_dqdPE5) enable((*inhigh*) EN_dtau_vec_in_R7_dqdPE5) ;
    method dtau_vec_in_R1_dqdPE6(dtau_vec_in_R1_dqdPE6) enable((*inhigh*) EN_dtau_vec_in_R1_dqdPE6) ;
    method dtau_vec_in_R2_dqdPE6(dtau_vec_in_R2_dqdPE6) enable((*inhigh*) EN_dtau_vec_in_R2_dqdPE6) ;
    method dtau_vec_in_R3_dqdPE6(dtau_vec_in_R3_dqdPE6) enable((*inhigh*) EN_dtau_vec_in_R3_dqdPE6) ;
    method dtau_vec_in_R4_dqdPE6(dtau_vec_in_R4_dqdPE6) enable((*inhigh*) EN_dtau_vec_in_R4_dqdPE6) ;
    method dtau_vec_in_R5_dqdPE6(dtau_vec_in_R5_dqdPE6) enable((*inhigh*) EN_dtau_vec_in_R5_dqdPE6) ;
    method dtau_vec_in_R6_dqdPE6(dtau_vec_in_R6_dqdPE6) enable((*inhigh*) EN_dtau_vec_in_R6_dqdPE6) ;
    method dtau_vec_in_R7_dqdPE6(dtau_vec_in_R7_dqdPE6) enable((*inhigh*) EN_dtau_vec_in_R7_dqdPE6) ;
    method dtau_vec_in_R1_dqdPE7(dtau_vec_in_R1_dqdPE7) enable((*inhigh*) EN_dtau_vec_in_R1_dqdPE7) ;
    method dtau_vec_in_R2_dqdPE7(dtau_vec_in_R2_dqdPE7) enable((*inhigh*) EN_dtau_vec_in_R2_dqdPE7) ;
    method dtau_vec_in_R3_dqdPE7(dtau_vec_in_R3_dqdPE7) enable((*inhigh*) EN_dtau_vec_in_R3_dqdPE7) ;
    method dtau_vec_in_R4_dqdPE7(dtau_vec_in_R4_dqdPE7) enable((*inhigh*) EN_dtau_vec_in_R4_dqdPE7) ;
    method dtau_vec_in_R5_dqdPE7(dtau_vec_in_R5_dqdPE7) enable((*inhigh*) EN_dtau_vec_in_R5_dqdPE7) ;
    method dtau_vec_in_R6_dqdPE7(dtau_vec_in_R6_dqdPE7) enable((*inhigh*) EN_dtau_vec_in_R6_dqdPE7) ;
    method dtau_vec_in_R7_dqdPE7(dtau_vec_in_R7_dqdPE7) enable((*inhigh*) EN_dtau_vec_in_R7_dqdPE7) ;

    method output_ready output_ready();
    method output_ready_minv output_ready_minv();
    method tau_curr_out_rnea tau_curr_out_rnea();


    method f_upd_prev_vec_out_AX_rnea f_upd_prev_vec_out_AX_rnea();
    method f_upd_prev_vec_out_AY_rnea f_upd_prev_vec_out_AY_rnea();
    method f_upd_prev_vec_out_AZ_rnea f_upd_prev_vec_out_AZ_rnea();
    method f_upd_prev_vec_out_LX_rnea f_upd_prev_vec_out_LX_rnea();
    method f_upd_prev_vec_out_LY_rnea f_upd_prev_vec_out_LY_rnea();
    method f_upd_prev_vec_out_LZ_rnea f_upd_prev_vec_out_LZ_rnea();

    method dtau_curr_out_dqPE1 dtau_curr_out_dqPE1();
    method dtau_curr_out_dqPE2 dtau_curr_out_dqPE2();
    method dtau_curr_out_dqPE3 dtau_curr_out_dqPE3();
    method dtau_curr_out_dqPE4 dtau_curr_out_dqPE4();
    method dtau_curr_out_dqPE5 dtau_curr_out_dqPE5();
    method dtau_curr_out_dqPE6 dtau_curr_out_dqPE6();
    method dtau_curr_out_dqPE7 dtau_curr_out_dqPE7();
    method dtau_curr_out_dqdPE1 dtau_curr_out_dqdPE1();
    method dtau_curr_out_dqdPE2 dtau_curr_out_dqdPE2();
    method dtau_curr_out_dqdPE3 dtau_curr_out_dqdPE3();
    method dtau_curr_out_dqdPE4 dtau_curr_out_dqdPE4();
    method dtau_curr_out_dqdPE5 dtau_curr_out_dqdPE5();
    method dtau_curr_out_dqdPE6 dtau_curr_out_dqdPE6();
    method dtau_curr_out_dqdPE7 dtau_curr_out_dqdPE7();
    method dfdq_upd_prev_vec_out_AX_dqPE1 dfdq_upd_prev_vec_out_AX_dqPE1();
    method dfdq_upd_prev_vec_out_AY_dqPE1 dfdq_upd_prev_vec_out_AY_dqPE1();
    method dfdq_upd_prev_vec_out_AZ_dqPE1 dfdq_upd_prev_vec_out_AZ_dqPE1();
    method dfdq_upd_prev_vec_out_LX_dqPE1 dfdq_upd_prev_vec_out_LX_dqPE1();
    method dfdq_upd_prev_vec_out_LY_dqPE1 dfdq_upd_prev_vec_out_LY_dqPE1();
    method dfdq_upd_prev_vec_out_LZ_dqPE1 dfdq_upd_prev_vec_out_LZ_dqPE1();
    method dfdq_upd_prev_vec_out_AX_dqPE2 dfdq_upd_prev_vec_out_AX_dqPE2();
    method dfdq_upd_prev_vec_out_AY_dqPE2 dfdq_upd_prev_vec_out_AY_dqPE2();
    method dfdq_upd_prev_vec_out_AZ_dqPE2 dfdq_upd_prev_vec_out_AZ_dqPE2();
    method dfdq_upd_prev_vec_out_LX_dqPE2 dfdq_upd_prev_vec_out_LX_dqPE2();
    method dfdq_upd_prev_vec_out_LY_dqPE2 dfdq_upd_prev_vec_out_LY_dqPE2();
    method dfdq_upd_prev_vec_out_LZ_dqPE2 dfdq_upd_prev_vec_out_LZ_dqPE2();
    method dfdq_upd_prev_vec_out_AX_dqPE3 dfdq_upd_prev_vec_out_AX_dqPE3();
    method dfdq_upd_prev_vec_out_AY_dqPE3 dfdq_upd_prev_vec_out_AY_dqPE3();
    method dfdq_upd_prev_vec_out_AZ_dqPE3 dfdq_upd_prev_vec_out_AZ_dqPE3();
    method dfdq_upd_prev_vec_out_LX_dqPE3 dfdq_upd_prev_vec_out_LX_dqPE3();
    method dfdq_upd_prev_vec_out_LY_dqPE3 dfdq_upd_prev_vec_out_LY_dqPE3();
    method dfdq_upd_prev_vec_out_LZ_dqPE3 dfdq_upd_prev_vec_out_LZ_dqPE3();
    method dfdq_upd_prev_vec_out_AX_dqPE4 dfdq_upd_prev_vec_out_AX_dqPE4();
    method dfdq_upd_prev_vec_out_AY_dqPE4 dfdq_upd_prev_vec_out_AY_dqPE4();
    method dfdq_upd_prev_vec_out_AZ_dqPE4 dfdq_upd_prev_vec_out_AZ_dqPE4();
    method dfdq_upd_prev_vec_out_LX_dqPE4 dfdq_upd_prev_vec_out_LX_dqPE4();
    method dfdq_upd_prev_vec_out_LY_dqPE4 dfdq_upd_prev_vec_out_LY_dqPE4();
    method dfdq_upd_prev_vec_out_LZ_dqPE4 dfdq_upd_prev_vec_out_LZ_dqPE4();
    method dfdq_upd_prev_vec_out_AX_dqPE5 dfdq_upd_prev_vec_out_AX_dqPE5();
    method dfdq_upd_prev_vec_out_AY_dqPE5 dfdq_upd_prev_vec_out_AY_dqPE5();
    method dfdq_upd_prev_vec_out_AZ_dqPE5 dfdq_upd_prev_vec_out_AZ_dqPE5();
    method dfdq_upd_prev_vec_out_LX_dqPE5 dfdq_upd_prev_vec_out_LX_dqPE5();
    method dfdq_upd_prev_vec_out_LY_dqPE5 dfdq_upd_prev_vec_out_LY_dqPE5();
    method dfdq_upd_prev_vec_out_LZ_dqPE5 dfdq_upd_prev_vec_out_LZ_dqPE5();
    method dfdq_upd_prev_vec_out_AX_dqPE6 dfdq_upd_prev_vec_out_AX_dqPE6();
    method dfdq_upd_prev_vec_out_AY_dqPE6 dfdq_upd_prev_vec_out_AY_dqPE6();
    method dfdq_upd_prev_vec_out_AZ_dqPE6 dfdq_upd_prev_vec_out_AZ_dqPE6();
    method dfdq_upd_prev_vec_out_LX_dqPE6 dfdq_upd_prev_vec_out_LX_dqPE6();
    method dfdq_upd_prev_vec_out_LY_dqPE6 dfdq_upd_prev_vec_out_LY_dqPE6();
    method dfdq_upd_prev_vec_out_LZ_dqPE6 dfdq_upd_prev_vec_out_LZ_dqPE6();
    method dfdq_upd_prev_vec_out_AX_dqPE7 dfdq_upd_prev_vec_out_AX_dqPE7();
    method dfdq_upd_prev_vec_out_AY_dqPE7 dfdq_upd_prev_vec_out_AY_dqPE7();
    method dfdq_upd_prev_vec_out_AZ_dqPE7 dfdq_upd_prev_vec_out_AZ_dqPE7();
    method dfdq_upd_prev_vec_out_LX_dqPE7 dfdq_upd_prev_vec_out_LX_dqPE7();
    method dfdq_upd_prev_vec_out_LY_dqPE7 dfdq_upd_prev_vec_out_LY_dqPE7();
    method dfdq_upd_prev_vec_out_LZ_dqPE7 dfdq_upd_prev_vec_out_LZ_dqPE7();
    method dfdqd_upd_prev_vec_out_AX_dqdPE1 dfdqd_upd_prev_vec_out_AX_dqdPE1();
    method dfdqd_upd_prev_vec_out_AY_dqdPE1 dfdqd_upd_prev_vec_out_AY_dqdPE1();
    method dfdqd_upd_prev_vec_out_AZ_dqdPE1 dfdqd_upd_prev_vec_out_AZ_dqdPE1();
    method dfdqd_upd_prev_vec_out_LX_dqdPE1 dfdqd_upd_prev_vec_out_LX_dqdPE1();
    method dfdqd_upd_prev_vec_out_LY_dqdPE1 dfdqd_upd_prev_vec_out_LY_dqdPE1();
    method dfdqd_upd_prev_vec_out_LZ_dqdPE1 dfdqd_upd_prev_vec_out_LZ_dqdPE1();
    method dfdqd_upd_prev_vec_out_AX_dqdPE2 dfdqd_upd_prev_vec_out_AX_dqdPE2();
    method dfdqd_upd_prev_vec_out_AY_dqdPE2 dfdqd_upd_prev_vec_out_AY_dqdPE2();
    method dfdqd_upd_prev_vec_out_AZ_dqdPE2 dfdqd_upd_prev_vec_out_AZ_dqdPE2();
    method dfdqd_upd_prev_vec_out_LX_dqdPE2 dfdqd_upd_prev_vec_out_LX_dqdPE2();
    method dfdqd_upd_prev_vec_out_LY_dqdPE2 dfdqd_upd_prev_vec_out_LY_dqdPE2();
    method dfdqd_upd_prev_vec_out_LZ_dqdPE2 dfdqd_upd_prev_vec_out_LZ_dqdPE2();
    method dfdqd_upd_prev_vec_out_AX_dqdPE3 dfdqd_upd_prev_vec_out_AX_dqdPE3();
    method dfdqd_upd_prev_vec_out_AY_dqdPE3 dfdqd_upd_prev_vec_out_AY_dqdPE3();
    method dfdqd_upd_prev_vec_out_AZ_dqdPE3 dfdqd_upd_prev_vec_out_AZ_dqdPE3();
    method dfdqd_upd_prev_vec_out_LX_dqdPE3 dfdqd_upd_prev_vec_out_LX_dqdPE3();
    method dfdqd_upd_prev_vec_out_LY_dqdPE3 dfdqd_upd_prev_vec_out_LY_dqdPE3();
    method dfdqd_upd_prev_vec_out_LZ_dqdPE3 dfdqd_upd_prev_vec_out_LZ_dqdPE3();
    method dfdqd_upd_prev_vec_out_AX_dqdPE4 dfdqd_upd_prev_vec_out_AX_dqdPE4();
    method dfdqd_upd_prev_vec_out_AY_dqdPE4 dfdqd_upd_prev_vec_out_AY_dqdPE4();
    method dfdqd_upd_prev_vec_out_AZ_dqdPE4 dfdqd_upd_prev_vec_out_AZ_dqdPE4();
    method dfdqd_upd_prev_vec_out_LX_dqdPE4 dfdqd_upd_prev_vec_out_LX_dqdPE4();
    method dfdqd_upd_prev_vec_out_LY_dqdPE4 dfdqd_upd_prev_vec_out_LY_dqdPE4();
    method dfdqd_upd_prev_vec_out_LZ_dqdPE4 dfdqd_upd_prev_vec_out_LZ_dqdPE4();
    method dfdqd_upd_prev_vec_out_AX_dqdPE5 dfdqd_upd_prev_vec_out_AX_dqdPE5();
    method dfdqd_upd_prev_vec_out_AY_dqdPE5 dfdqd_upd_prev_vec_out_AY_dqdPE5();
    method dfdqd_upd_prev_vec_out_AZ_dqdPE5 dfdqd_upd_prev_vec_out_AZ_dqdPE5();
    method dfdqd_upd_prev_vec_out_LX_dqdPE5 dfdqd_upd_prev_vec_out_LX_dqdPE5();
    method dfdqd_upd_prev_vec_out_LY_dqdPE5 dfdqd_upd_prev_vec_out_LY_dqdPE5();
    method dfdqd_upd_prev_vec_out_LZ_dqdPE5 dfdqd_upd_prev_vec_out_LZ_dqdPE5();
    method dfdqd_upd_prev_vec_out_AX_dqdPE6 dfdqd_upd_prev_vec_out_AX_dqdPE6();
    method dfdqd_upd_prev_vec_out_AY_dqdPE6 dfdqd_upd_prev_vec_out_AY_dqdPE6();
    method dfdqd_upd_prev_vec_out_AZ_dqdPE6 dfdqd_upd_prev_vec_out_AZ_dqdPE6();
    method dfdqd_upd_prev_vec_out_LX_dqdPE6 dfdqd_upd_prev_vec_out_LX_dqdPE6();
    method dfdqd_upd_prev_vec_out_LY_dqdPE6 dfdqd_upd_prev_vec_out_LY_dqdPE6();
    method dfdqd_upd_prev_vec_out_LZ_dqdPE6 dfdqd_upd_prev_vec_out_LZ_dqdPE6();
    method dfdqd_upd_prev_vec_out_AX_dqdPE7 dfdqd_upd_prev_vec_out_AX_dqdPE7();
    method dfdqd_upd_prev_vec_out_AY_dqdPE7 dfdqd_upd_prev_vec_out_AY_dqdPE7();
    method dfdqd_upd_prev_vec_out_AZ_dqdPE7 dfdqd_upd_prev_vec_out_AZ_dqdPE7();
    method dfdqd_upd_prev_vec_out_LX_dqdPE7 dfdqd_upd_prev_vec_out_LX_dqdPE7();
    method dfdqd_upd_prev_vec_out_LY_dqdPE7 dfdqd_upd_prev_vec_out_LY_dqdPE7();
    method dfdqd_upd_prev_vec_out_LZ_dqdPE7 dfdqd_upd_prev_vec_out_LZ_dqdPE7();
    method minv_vec_out_R1_dqdPE1 minv_vec_out_R1_dqdPE1();
    method minv_vec_out_R2_dqdPE1 minv_vec_out_R2_dqdPE1();
    method minv_vec_out_R3_dqdPE1 minv_vec_out_R3_dqdPE1();
    method minv_vec_out_R4_dqdPE1 minv_vec_out_R4_dqdPE1();
    method minv_vec_out_R5_dqdPE1 minv_vec_out_R5_dqdPE1();
    method minv_vec_out_R6_dqdPE1 minv_vec_out_R6_dqdPE1();
    method minv_vec_out_R7_dqdPE1 minv_vec_out_R7_dqdPE1();
    method minv_vec_out_R1_dqdPE2 minv_vec_out_R1_dqdPE2();
    method minv_vec_out_R2_dqdPE2 minv_vec_out_R2_dqdPE2();
    method minv_vec_out_R3_dqdPE2 minv_vec_out_R3_dqdPE2();
    method minv_vec_out_R4_dqdPE2 minv_vec_out_R4_dqdPE2();
    method minv_vec_out_R5_dqdPE2 minv_vec_out_R5_dqdPE2();
    method minv_vec_out_R6_dqdPE2 minv_vec_out_R6_dqdPE2();
    method minv_vec_out_R7_dqdPE2 minv_vec_out_R7_dqdPE2();
    method minv_vec_out_R1_dqdPE3 minv_vec_out_R1_dqdPE3();
    method minv_vec_out_R2_dqdPE3 minv_vec_out_R2_dqdPE3();
    method minv_vec_out_R3_dqdPE3 minv_vec_out_R3_dqdPE3();
    method minv_vec_out_R4_dqdPE3 minv_vec_out_R4_dqdPE3();
    method minv_vec_out_R5_dqdPE3 minv_vec_out_R5_dqdPE3();
    method minv_vec_out_R6_dqdPE3 minv_vec_out_R6_dqdPE3();
    method minv_vec_out_R7_dqdPE3 minv_vec_out_R7_dqdPE3();
    method minv_vec_out_R1_dqdPE4 minv_vec_out_R1_dqdPE4();
    method minv_vec_out_R2_dqdPE4 minv_vec_out_R2_dqdPE4();
    method minv_vec_out_R3_dqdPE4 minv_vec_out_R3_dqdPE4();
    method minv_vec_out_R4_dqdPE4 minv_vec_out_R4_dqdPE4();
    method minv_vec_out_R5_dqdPE4 minv_vec_out_R5_dqdPE4();
    method minv_vec_out_R6_dqdPE4 minv_vec_out_R6_dqdPE4();
    method minv_vec_out_R7_dqdPE4 minv_vec_out_R7_dqdPE4();
    method minv_vec_out_R1_dqdPE5 minv_vec_out_R1_dqdPE5();
    method minv_vec_out_R2_dqdPE5 minv_vec_out_R2_dqdPE5();
    method minv_vec_out_R3_dqdPE5 minv_vec_out_R3_dqdPE5();
    method minv_vec_out_R4_dqdPE5 minv_vec_out_R4_dqdPE5();
    method minv_vec_out_R5_dqdPE5 minv_vec_out_R5_dqdPE5();
    method minv_vec_out_R6_dqdPE5 minv_vec_out_R6_dqdPE5();
    method minv_vec_out_R7_dqdPE5 minv_vec_out_R7_dqdPE5();
    method minv_vec_out_R1_dqdPE6 minv_vec_out_R1_dqdPE6();
    method minv_vec_out_R2_dqdPE6 minv_vec_out_R2_dqdPE6();
    method minv_vec_out_R3_dqdPE6 minv_vec_out_R3_dqdPE6();
    method minv_vec_out_R4_dqdPE6 minv_vec_out_R4_dqdPE6();
    method minv_vec_out_R5_dqdPE6 minv_vec_out_R5_dqdPE6();
    method minv_vec_out_R6_dqdPE6 minv_vec_out_R6_dqdPE6();
    method minv_vec_out_R7_dqdPE6 minv_vec_out_R7_dqdPE6();
    method minv_vec_out_R1_dqdPE7 minv_vec_out_R1_dqdPE7();
    method minv_vec_out_R2_dqdPE7 minv_vec_out_R2_dqdPE7();
    method minv_vec_out_R3_dqdPE7 minv_vec_out_R3_dqdPE7();
    method minv_vec_out_R4_dqdPE7 minv_vec_out_R4_dqdPE7();
    method minv_vec_out_R5_dqdPE7 minv_vec_out_R5_dqdPE7();
    method minv_vec_out_R6_dqdPE7 minv_vec_out_R6_dqdPE7();
    method minv_vec_out_R7_dqdPE7 minv_vec_out_R7_dqdPE7();

    schedule (
        get_data, get_data_minv, link_in_rnea, sinq_val_in_rnea, cosq_val_in_rnea,
        f_upd_curr_vec_in_AX_rnea, f_upd_curr_vec_in_AY_rnea, f_upd_curr_vec_in_AZ_rnea, f_upd_curr_vec_in_LX_rnea, f_upd_curr_vec_in_LY_rnea, f_upd_curr_vec_in_LZ_rnea, f_prev_vec_in_AX_rnea, f_prev_vec_in_AY_rnea, f_prev_vec_in_AZ_rnea, f_prev_vec_in_LX_rnea, f_prev_vec_in_LY_rnea, f_prev_vec_in_LZ_rnea,
        link_in_dqPE1, link_in_dqPE2, link_in_dqPE3, link_in_dqPE4, link_in_dqPE5, link_in_dqPE6, link_in_dqPE7, link_in_dqdPE1, link_in_dqdPE2, link_in_dqdPE3, link_in_dqdPE4, link_in_dqdPE5, link_in_dqdPE6, link_in_dqdPE7, derv_in_dqPE1, derv_in_dqPE2, derv_in_dqPE3, derv_in_dqPE4, derv_in_dqPE5, derv_in_dqPE6, derv_in_dqPE7, derv_in_dqdPE1, derv_in_dqdPE2, derv_in_dqdPE3, derv_in_dqdPE4, derv_in_dqdPE5, derv_in_dqdPE6, derv_in_dqdPE7,
        sinq_val_in_dqPE1, sinq_val_in_dqPE2, sinq_val_in_dqPE3, sinq_val_in_dqPE4, sinq_val_in_dqPE5, sinq_val_in_dqPE6, sinq_val_in_dqPE7, sinq_val_in_dqdPE1, sinq_val_in_dqdPE2, sinq_val_in_dqdPE3, sinq_val_in_dqdPE4, sinq_val_in_dqdPE5, sinq_val_in_dqdPE6, sinq_val_in_dqdPE7, cosq_val_in_dqPE1, cosq_val_in_dqPE2, cosq_val_in_dqPE3, cosq_val_in_dqPE4, cosq_val_in_dqPE5, cosq_val_in_dqPE6, cosq_val_in_dqPE7, cosq_val_in_dqdPE1, cosq_val_in_dqdPE2, cosq_val_in_dqdPE3, cosq_val_in_dqdPE4, cosq_val_in_dqdPE5, cosq_val_in_dqdPE6, cosq_val_in_dqdPE7,
        f_upd_curr_vec_in_AX_dqPE1, f_upd_curr_vec_in_AY_dqPE1, f_upd_curr_vec_in_AZ_dqPE1, f_upd_curr_vec_in_LX_dqPE1, f_upd_curr_vec_in_LY_dqPE1, f_upd_curr_vec_in_LZ_dqPE1, f_upd_curr_vec_in_AX_dqPE2, f_upd_curr_vec_in_AY_dqPE2, f_upd_curr_vec_in_AZ_dqPE2, f_upd_curr_vec_in_LX_dqPE2, f_upd_curr_vec_in_LY_dqPE2, f_upd_curr_vec_in_LZ_dqPE2, f_upd_curr_vec_in_AX_dqPE3, f_upd_curr_vec_in_AY_dqPE3, f_upd_curr_vec_in_AZ_dqPE3, f_upd_curr_vec_in_LX_dqPE3, f_upd_curr_vec_in_LY_dqPE3, f_upd_curr_vec_in_LZ_dqPE3, f_upd_curr_vec_in_AX_dqPE4, f_upd_curr_vec_in_AY_dqPE4, f_upd_curr_vec_in_AZ_dqPE4, f_upd_curr_vec_in_LX_dqPE4, f_upd_curr_vec_in_LY_dqPE4, f_upd_curr_vec_in_LZ_dqPE4, f_upd_curr_vec_in_AX_dqPE5, f_upd_curr_vec_in_AY_dqPE5, f_upd_curr_vec_in_AZ_dqPE5, f_upd_curr_vec_in_LX_dqPE5, f_upd_curr_vec_in_LY_dqPE5, f_upd_curr_vec_in_LZ_dqPE5, f_upd_curr_vec_in_AX_dqPE6, f_upd_curr_vec_in_AY_dqPE6, f_upd_curr_vec_in_AZ_dqPE6, f_upd_curr_vec_in_LX_dqPE6, f_upd_curr_vec_in_LY_dqPE6, f_upd_curr_vec_in_LZ_dqPE6, f_upd_curr_vec_in_AX_dqPE7, f_upd_curr_vec_in_AY_dqPE7, f_upd_curr_vec_in_AZ_dqPE7, f_upd_curr_vec_in_LX_dqPE7, f_upd_curr_vec_in_LY_dqPE7, f_upd_curr_vec_in_LZ_dqPE7, dfdq_prev_vec_in_AX_dqPE1, dfdq_prev_vec_in_AY_dqPE1, dfdq_prev_vec_in_AZ_dqPE1, dfdq_prev_vec_in_LX_dqPE1, dfdq_prev_vec_in_LY_dqPE1, dfdq_prev_vec_in_LZ_dqPE1, dfdq_prev_vec_in_AX_dqPE2, dfdq_prev_vec_in_AY_dqPE2, dfdq_prev_vec_in_AZ_dqPE2, dfdq_prev_vec_in_LX_dqPE2, dfdq_prev_vec_in_LY_dqPE2, dfdq_prev_vec_in_LZ_dqPE2, dfdq_prev_vec_in_AX_dqPE3, dfdq_prev_vec_in_AY_dqPE3, dfdq_prev_vec_in_AZ_dqPE3, dfdq_prev_vec_in_LX_dqPE3, dfdq_prev_vec_in_LY_dqPE3, dfdq_prev_vec_in_LZ_dqPE3, dfdq_prev_vec_in_AX_dqPE4, dfdq_prev_vec_in_AY_dqPE4, dfdq_prev_vec_in_AZ_dqPE4, dfdq_prev_vec_in_LX_dqPE4, dfdq_prev_vec_in_LY_dqPE4, dfdq_prev_vec_in_LZ_dqPE4, dfdq_prev_vec_in_AX_dqPE5, dfdq_prev_vec_in_AY_dqPE5, dfdq_prev_vec_in_AZ_dqPE5, dfdq_prev_vec_in_LX_dqPE5, dfdq_prev_vec_in_LY_dqPE5, dfdq_prev_vec_in_LZ_dqPE5, dfdq_prev_vec_in_AX_dqPE6, dfdq_prev_vec_in_AY_dqPE6, dfdq_prev_vec_in_AZ_dqPE6, dfdq_prev_vec_in_LX_dqPE6, dfdq_prev_vec_in_LY_dqPE6, dfdq_prev_vec_in_LZ_dqPE6, dfdq_prev_vec_in_AX_dqPE7, dfdq_prev_vec_in_AY_dqPE7, dfdq_prev_vec_in_AZ_dqPE7, dfdq_prev_vec_in_LX_dqPE7, dfdq_prev_vec_in_LY_dqPE7, dfdq_prev_vec_in_LZ_dqPE7, dfdq_upd_curr_vec_in_AX_dqPE1, dfdq_upd_curr_vec_in_AY_dqPE1, dfdq_upd_curr_vec_in_AZ_dqPE1, dfdq_upd_curr_vec_in_LX_dqPE1, dfdq_upd_curr_vec_in_LY_dqPE1, dfdq_upd_curr_vec_in_LZ_dqPE1, dfdq_upd_curr_vec_in_AX_dqPE2, dfdq_upd_curr_vec_in_AY_dqPE2, dfdq_upd_curr_vec_in_AZ_dqPE2, dfdq_upd_curr_vec_in_LX_dqPE2, dfdq_upd_curr_vec_in_LY_dqPE2, dfdq_upd_curr_vec_in_LZ_dqPE2, dfdq_upd_curr_vec_in_AX_dqPE3, dfdq_upd_curr_vec_in_AY_dqPE3, dfdq_upd_curr_vec_in_AZ_dqPE3, dfdq_upd_curr_vec_in_LX_dqPE3, dfdq_upd_curr_vec_in_LY_dqPE3, dfdq_upd_curr_vec_in_LZ_dqPE3, dfdq_upd_curr_vec_in_AX_dqPE4, dfdq_upd_curr_vec_in_AY_dqPE4, dfdq_upd_curr_vec_in_AZ_dqPE4, dfdq_upd_curr_vec_in_LX_dqPE4, dfdq_upd_curr_vec_in_LY_dqPE4, dfdq_upd_curr_vec_in_LZ_dqPE4, dfdq_upd_curr_vec_in_AX_dqPE5, dfdq_upd_curr_vec_in_AY_dqPE5, dfdq_upd_curr_vec_in_AZ_dqPE5, dfdq_upd_curr_vec_in_LX_dqPE5, dfdq_upd_curr_vec_in_LY_dqPE5, dfdq_upd_curr_vec_in_LZ_dqPE5, dfdq_upd_curr_vec_in_AX_dqPE6, dfdq_upd_curr_vec_in_AY_dqPE6, dfdq_upd_curr_vec_in_AZ_dqPE6, dfdq_upd_curr_vec_in_LX_dqPE6, dfdq_upd_curr_vec_in_LY_dqPE6, dfdq_upd_curr_vec_in_LZ_dqPE6, dfdq_upd_curr_vec_in_AX_dqPE7, dfdq_upd_curr_vec_in_AY_dqPE7, dfdq_upd_curr_vec_in_AZ_dqPE7, dfdq_upd_curr_vec_in_LX_dqPE7, dfdq_upd_curr_vec_in_LY_dqPE7, dfdq_upd_curr_vec_in_LZ_dqPE7, dfdqd_prev_vec_in_AX_dqdPE1, dfdqd_prev_vec_in_AY_dqdPE1, dfdqd_prev_vec_in_AZ_dqdPE1, dfdqd_prev_vec_in_LX_dqdPE1, dfdqd_prev_vec_in_LY_dqdPE1, dfdqd_prev_vec_in_LZ_dqdPE1, dfdqd_prev_vec_in_AX_dqdPE2, dfdqd_prev_vec_in_AY_dqdPE2, dfdqd_prev_vec_in_AZ_dqdPE2, dfdqd_prev_vec_in_LX_dqdPE2, dfdqd_prev_vec_in_LY_dqdPE2, dfdqd_prev_vec_in_LZ_dqdPE2, dfdqd_prev_vec_in_AX_dqdPE3, dfdqd_prev_vec_in_AY_dqdPE3, dfdqd_prev_vec_in_AZ_dqdPE3, dfdqd_prev_vec_in_LX_dqdPE3, dfdqd_prev_vec_in_LY_dqdPE3, dfdqd_prev_vec_in_LZ_dqdPE3, dfdqd_prev_vec_in_AX_dqdPE4, dfdqd_prev_vec_in_AY_dqdPE4, dfdqd_prev_vec_in_AZ_dqdPE4, dfdqd_prev_vec_in_LX_dqdPE4, dfdqd_prev_vec_in_LY_dqdPE4, dfdqd_prev_vec_in_LZ_dqdPE4, dfdqd_prev_vec_in_AX_dqdPE5, dfdqd_prev_vec_in_AY_dqdPE5, dfdqd_prev_vec_in_AZ_dqdPE5, dfdqd_prev_vec_in_LX_dqdPE5, dfdqd_prev_vec_in_LY_dqdPE5, dfdqd_prev_vec_in_LZ_dqdPE5, dfdqd_prev_vec_in_AX_dqdPE6, dfdqd_prev_vec_in_AY_dqdPE6, dfdqd_prev_vec_in_AZ_dqdPE6, dfdqd_prev_vec_in_LX_dqdPE6, dfdqd_prev_vec_in_LY_dqdPE6, dfdqd_prev_vec_in_LZ_dqdPE6, dfdqd_prev_vec_in_AX_dqdPE7, dfdqd_prev_vec_in_AY_dqdPE7, dfdqd_prev_vec_in_AZ_dqdPE7, dfdqd_prev_vec_in_LX_dqdPE7, dfdqd_prev_vec_in_LY_dqdPE7, dfdqd_prev_vec_in_LZ_dqdPE7, dfdqd_upd_curr_vec_in_AX_dqdPE1, dfdqd_upd_curr_vec_in_AY_dqdPE1, dfdqd_upd_curr_vec_in_AZ_dqdPE1, dfdqd_upd_curr_vec_in_LX_dqdPE1, dfdqd_upd_curr_vec_in_LY_dqdPE1, dfdqd_upd_curr_vec_in_LZ_dqdPE1, dfdqd_upd_curr_vec_in_AX_dqdPE2, dfdqd_upd_curr_vec_in_AY_dqdPE2, dfdqd_upd_curr_vec_in_AZ_dqdPE2, dfdqd_upd_curr_vec_in_LX_dqdPE2, dfdqd_upd_curr_vec_in_LY_dqdPE2, dfdqd_upd_curr_vec_in_LZ_dqdPE2, dfdqd_upd_curr_vec_in_AX_dqdPE3, dfdqd_upd_curr_vec_in_AY_dqdPE3, dfdqd_upd_curr_vec_in_AZ_dqdPE3, dfdqd_upd_curr_vec_in_LX_dqdPE3, dfdqd_upd_curr_vec_in_LY_dqdPE3, dfdqd_upd_curr_vec_in_LZ_dqdPE3, dfdqd_upd_curr_vec_in_AX_dqdPE4, dfdqd_upd_curr_vec_in_AY_dqdPE4, dfdqd_upd_curr_vec_in_AZ_dqdPE4, dfdqd_upd_curr_vec_in_LX_dqdPE4, dfdqd_upd_curr_vec_in_LY_dqdPE4, dfdqd_upd_curr_vec_in_LZ_dqdPE4, dfdqd_upd_curr_vec_in_AX_dqdPE5, dfdqd_upd_curr_vec_in_AY_dqdPE5, dfdqd_upd_curr_vec_in_AZ_dqdPE5, dfdqd_upd_curr_vec_in_LX_dqdPE5, dfdqd_upd_curr_vec_in_LY_dqdPE5, dfdqd_upd_curr_vec_in_LZ_dqdPE5, dfdqd_upd_curr_vec_in_AX_dqdPE6, dfdqd_upd_curr_vec_in_AY_dqdPE6, dfdqd_upd_curr_vec_in_AZ_dqdPE6, dfdqd_upd_curr_vec_in_LX_dqdPE6, dfdqd_upd_curr_vec_in_LY_dqdPE6, dfdqd_upd_curr_vec_in_LZ_dqdPE6, dfdqd_upd_curr_vec_in_AX_dqdPE7, dfdqd_upd_curr_vec_in_AY_dqdPE7, dfdqd_upd_curr_vec_in_AZ_dqdPE7, dfdqd_upd_curr_vec_in_LX_dqdPE7, dfdqd_upd_curr_vec_in_LY_dqdPE7, dfdqd_upd_curr_vec_in_LZ_dqdPE7,
        minv_block_in_R1_C1_dqdPE1, minv_block_in_R2_C1_dqdPE1, minv_block_in_R3_C1_dqdPE1, minv_block_in_R4_C1_dqdPE1, minv_block_in_R5_C1_dqdPE1, minv_block_in_R6_C1_dqdPE1, minv_block_in_R7_C1_dqdPE1, minv_block_in_R1_C2_dqdPE1, minv_block_in_R2_C2_dqdPE1, minv_block_in_R3_C2_dqdPE1, minv_block_in_R4_C2_dqdPE1, minv_block_in_R5_C2_dqdPE1, minv_block_in_R6_C2_dqdPE1, minv_block_in_R7_C2_dqdPE1, minv_block_in_R1_C3_dqdPE1, minv_block_in_R2_C3_dqdPE1, minv_block_in_R3_C3_dqdPE1, minv_block_in_R4_C3_dqdPE1, minv_block_in_R5_C3_dqdPE1, minv_block_in_R6_C3_dqdPE1, minv_block_in_R7_C3_dqdPE1, minv_block_in_R1_C4_dqdPE1, minv_block_in_R2_C4_dqdPE1, minv_block_in_R3_C4_dqdPE1, minv_block_in_R4_C4_dqdPE1, minv_block_in_R5_C4_dqdPE1, minv_block_in_R6_C4_dqdPE1, minv_block_in_R7_C4_dqdPE1, minv_block_in_R1_C5_dqdPE1, minv_block_in_R2_C5_dqdPE1, minv_block_in_R3_C5_dqdPE1, minv_block_in_R4_C5_dqdPE1, minv_block_in_R5_C5_dqdPE1, minv_block_in_R6_C5_dqdPE1, minv_block_in_R7_C5_dqdPE1, minv_block_in_R1_C6_dqdPE1, minv_block_in_R2_C6_dqdPE1, minv_block_in_R3_C6_dqdPE1, minv_block_in_R4_C6_dqdPE1, minv_block_in_R5_C6_dqdPE1, minv_block_in_R6_C6_dqdPE1, minv_block_in_R7_C6_dqdPE1, minv_block_in_R1_C7_dqdPE1, minv_block_in_R2_C7_dqdPE1, minv_block_in_R3_C7_dqdPE1, minv_block_in_R4_C7_dqdPE1, minv_block_in_R5_C7_dqdPE1, minv_block_in_R6_C7_dqdPE1, minv_block_in_R7_C7_dqdPE1, minv_block_in_R1_C1_dqdPE2, minv_block_in_R2_C1_dqdPE2, minv_block_in_R3_C1_dqdPE2, minv_block_in_R4_C1_dqdPE2, minv_block_in_R5_C1_dqdPE2, minv_block_in_R6_C1_dqdPE2, minv_block_in_R7_C1_dqdPE2, minv_block_in_R1_C2_dqdPE2, minv_block_in_R2_C2_dqdPE2, minv_block_in_R3_C2_dqdPE2, minv_block_in_R4_C2_dqdPE2, minv_block_in_R5_C2_dqdPE2, minv_block_in_R6_C2_dqdPE2, minv_block_in_R7_C2_dqdPE2, minv_block_in_R1_C3_dqdPE2, minv_block_in_R2_C3_dqdPE2, minv_block_in_R3_C3_dqdPE2, minv_block_in_R4_C3_dqdPE2, minv_block_in_R5_C3_dqdPE2, minv_block_in_R6_C3_dqdPE2, minv_block_in_R7_C3_dqdPE2, minv_block_in_R1_C4_dqdPE2, minv_block_in_R2_C4_dqdPE2, minv_block_in_R3_C4_dqdPE2, minv_block_in_R4_C4_dqdPE2, minv_block_in_R5_C4_dqdPE2, minv_block_in_R6_C4_dqdPE2, minv_block_in_R7_C4_dqdPE2, minv_block_in_R1_C5_dqdPE2, minv_block_in_R2_C5_dqdPE2, minv_block_in_R3_C5_dqdPE2, minv_block_in_R4_C5_dqdPE2, minv_block_in_R5_C5_dqdPE2, minv_block_in_R6_C5_dqdPE2, minv_block_in_R7_C5_dqdPE2, minv_block_in_R1_C6_dqdPE2, minv_block_in_R2_C6_dqdPE2, minv_block_in_R3_C6_dqdPE2, minv_block_in_R4_C6_dqdPE2, minv_block_in_R5_C6_dqdPE2, minv_block_in_R6_C6_dqdPE2, minv_block_in_R7_C6_dqdPE2, minv_block_in_R1_C7_dqdPE2, minv_block_in_R2_C7_dqdPE2, minv_block_in_R3_C7_dqdPE2, minv_block_in_R4_C7_dqdPE2, minv_block_in_R5_C7_dqdPE2, minv_block_in_R6_C7_dqdPE2, minv_block_in_R7_C7_dqdPE2, minv_block_in_R1_C1_dqdPE3, minv_block_in_R2_C1_dqdPE3, minv_block_in_R3_C1_dqdPE3, minv_block_in_R4_C1_dqdPE3, minv_block_in_R5_C1_dqdPE3, minv_block_in_R6_C1_dqdPE3, minv_block_in_R7_C1_dqdPE3, minv_block_in_R1_C2_dqdPE3, minv_block_in_R2_C2_dqdPE3, minv_block_in_R3_C2_dqdPE3, minv_block_in_R4_C2_dqdPE3, minv_block_in_R5_C2_dqdPE3, minv_block_in_R6_C2_dqdPE3, minv_block_in_R7_C2_dqdPE3, minv_block_in_R1_C3_dqdPE3, minv_block_in_R2_C3_dqdPE3, minv_block_in_R3_C3_dqdPE3, minv_block_in_R4_C3_dqdPE3, minv_block_in_R5_C3_dqdPE3, minv_block_in_R6_C3_dqdPE3, minv_block_in_R7_C3_dqdPE3, minv_block_in_R1_C4_dqdPE3, minv_block_in_R2_C4_dqdPE3, minv_block_in_R3_C4_dqdPE3, minv_block_in_R4_C4_dqdPE3, minv_block_in_R5_C4_dqdPE3, minv_block_in_R6_C4_dqdPE3, minv_block_in_R7_C4_dqdPE3, minv_block_in_R1_C5_dqdPE3, minv_block_in_R2_C5_dqdPE3, minv_block_in_R3_C5_dqdPE3, minv_block_in_R4_C5_dqdPE3, minv_block_in_R5_C5_dqdPE3, minv_block_in_R6_C5_dqdPE3, minv_block_in_R7_C5_dqdPE3, minv_block_in_R1_C6_dqdPE3, minv_block_in_R2_C6_dqdPE3, minv_block_in_R3_C6_dqdPE3, minv_block_in_R4_C6_dqdPE3, minv_block_in_R5_C6_dqdPE3, minv_block_in_R6_C6_dqdPE3, minv_block_in_R7_C6_dqdPE3, minv_block_in_R1_C7_dqdPE3, minv_block_in_R2_C7_dqdPE3, minv_block_in_R3_C7_dqdPE3, minv_block_in_R4_C7_dqdPE3, minv_block_in_R5_C7_dqdPE3, minv_block_in_R6_C7_dqdPE3, minv_block_in_R7_C7_dqdPE3, minv_block_in_R1_C1_dqdPE4, minv_block_in_R2_C1_dqdPE4, minv_block_in_R3_C1_dqdPE4, minv_block_in_R4_C1_dqdPE4, minv_block_in_R5_C1_dqdPE4, minv_block_in_R6_C1_dqdPE4, minv_block_in_R7_C1_dqdPE4, minv_block_in_R1_C2_dqdPE4, minv_block_in_R2_C2_dqdPE4, minv_block_in_R3_C2_dqdPE4, minv_block_in_R4_C2_dqdPE4, minv_block_in_R5_C2_dqdPE4, minv_block_in_R6_C2_dqdPE4, minv_block_in_R7_C2_dqdPE4, minv_block_in_R1_C3_dqdPE4, minv_block_in_R2_C3_dqdPE4, minv_block_in_R3_C3_dqdPE4, minv_block_in_R4_C3_dqdPE4, minv_block_in_R5_C3_dqdPE4, minv_block_in_R6_C3_dqdPE4, minv_block_in_R7_C3_dqdPE4, minv_block_in_R1_C4_dqdPE4, minv_block_in_R2_C4_dqdPE4, minv_block_in_R3_C4_dqdPE4, minv_block_in_R4_C4_dqdPE4, minv_block_in_R5_C4_dqdPE4, minv_block_in_R6_C4_dqdPE4, minv_block_in_R7_C4_dqdPE4, minv_block_in_R1_C5_dqdPE4, minv_block_in_R2_C5_dqdPE4, minv_block_in_R3_C5_dqdPE4, minv_block_in_R4_C5_dqdPE4, minv_block_in_R5_C5_dqdPE4, minv_block_in_R6_C5_dqdPE4, minv_block_in_R7_C5_dqdPE4, minv_block_in_R1_C6_dqdPE4, minv_block_in_R2_C6_dqdPE4, minv_block_in_R3_C6_dqdPE4, minv_block_in_R4_C6_dqdPE4, minv_block_in_R5_C6_dqdPE4, minv_block_in_R6_C6_dqdPE4, minv_block_in_R7_C6_dqdPE4, minv_block_in_R1_C7_dqdPE4, minv_block_in_R2_C7_dqdPE4, minv_block_in_R3_C7_dqdPE4, minv_block_in_R4_C7_dqdPE4, minv_block_in_R5_C7_dqdPE4, minv_block_in_R6_C7_dqdPE4, minv_block_in_R7_C7_dqdPE4, minv_block_in_R1_C1_dqdPE5, minv_block_in_R2_C1_dqdPE5, minv_block_in_R3_C1_dqdPE5, minv_block_in_R4_C1_dqdPE5, minv_block_in_R5_C1_dqdPE5, minv_block_in_R6_C1_dqdPE5, minv_block_in_R7_C1_dqdPE5, minv_block_in_R1_C2_dqdPE5, minv_block_in_R2_C2_dqdPE5, minv_block_in_R3_C2_dqdPE5, minv_block_in_R4_C2_dqdPE5, minv_block_in_R5_C2_dqdPE5, minv_block_in_R6_C2_dqdPE5, minv_block_in_R7_C2_dqdPE5, minv_block_in_R1_C3_dqdPE5, minv_block_in_R2_C3_dqdPE5, minv_block_in_R3_C3_dqdPE5, minv_block_in_R4_C3_dqdPE5, minv_block_in_R5_C3_dqdPE5, minv_block_in_R6_C3_dqdPE5, minv_block_in_R7_C3_dqdPE5, minv_block_in_R1_C4_dqdPE5, minv_block_in_R2_C4_dqdPE5, minv_block_in_R3_C4_dqdPE5, minv_block_in_R4_C4_dqdPE5, minv_block_in_R5_C4_dqdPE5, minv_block_in_R6_C4_dqdPE5, minv_block_in_R7_C4_dqdPE5, minv_block_in_R1_C5_dqdPE5, minv_block_in_R2_C5_dqdPE5, minv_block_in_R3_C5_dqdPE5, minv_block_in_R4_C5_dqdPE5, minv_block_in_R5_C5_dqdPE5, minv_block_in_R6_C5_dqdPE5, minv_block_in_R7_C5_dqdPE5, minv_block_in_R1_C6_dqdPE5, minv_block_in_R2_C6_dqdPE5, minv_block_in_R3_C6_dqdPE5, minv_block_in_R4_C6_dqdPE5, minv_block_in_R5_C6_dqdPE5, minv_block_in_R6_C6_dqdPE5, minv_block_in_R7_C6_dqdPE5, minv_block_in_R1_C7_dqdPE5, minv_block_in_R2_C7_dqdPE5, minv_block_in_R3_C7_dqdPE5, minv_block_in_R4_C7_dqdPE5, minv_block_in_R5_C7_dqdPE5, minv_block_in_R6_C7_dqdPE5, minv_block_in_R7_C7_dqdPE5, minv_block_in_R1_C1_dqdPE6, minv_block_in_R2_C1_dqdPE6, minv_block_in_R3_C1_dqdPE6, minv_block_in_R4_C1_dqdPE6, minv_block_in_R5_C1_dqdPE6, minv_block_in_R6_C1_dqdPE6, minv_block_in_R7_C1_dqdPE6, minv_block_in_R1_C2_dqdPE6, minv_block_in_R2_C2_dqdPE6, minv_block_in_R3_C2_dqdPE6, minv_block_in_R4_C2_dqdPE6, minv_block_in_R5_C2_dqdPE6, minv_block_in_R6_C2_dqdPE6, minv_block_in_R7_C2_dqdPE6, minv_block_in_R1_C3_dqdPE6, minv_block_in_R2_C3_dqdPE6, minv_block_in_R3_C3_dqdPE6, minv_block_in_R4_C3_dqdPE6, minv_block_in_R5_C3_dqdPE6, minv_block_in_R6_C3_dqdPE6, minv_block_in_R7_C3_dqdPE6, minv_block_in_R1_C4_dqdPE6, minv_block_in_R2_C4_dqdPE6, minv_block_in_R3_C4_dqdPE6, minv_block_in_R4_C4_dqdPE6, minv_block_in_R5_C4_dqdPE6, minv_block_in_R6_C4_dqdPE6, minv_block_in_R7_C4_dqdPE6, minv_block_in_R1_C5_dqdPE6, minv_block_in_R2_C5_dqdPE6, minv_block_in_R3_C5_dqdPE6, minv_block_in_R4_C5_dqdPE6, minv_block_in_R5_C5_dqdPE6, minv_block_in_R6_C5_dqdPE6, minv_block_in_R7_C5_dqdPE6, minv_block_in_R1_C6_dqdPE6, minv_block_in_R2_C6_dqdPE6, minv_block_in_R3_C6_dqdPE6, minv_block_in_R4_C6_dqdPE6, minv_block_in_R5_C6_dqdPE6, minv_block_in_R6_C6_dqdPE6, minv_block_in_R7_C6_dqdPE6, minv_block_in_R1_C7_dqdPE6, minv_block_in_R2_C7_dqdPE6, minv_block_in_R3_C7_dqdPE6, minv_block_in_R4_C7_dqdPE6, minv_block_in_R5_C7_dqdPE6, minv_block_in_R6_C7_dqdPE6, minv_block_in_R7_C7_dqdPE6, minv_block_in_R1_C1_dqdPE7, minv_block_in_R2_C1_dqdPE7, minv_block_in_R3_C1_dqdPE7, minv_block_in_R4_C1_dqdPE7, minv_block_in_R5_C1_dqdPE7, minv_block_in_R6_C1_dqdPE7, minv_block_in_R7_C1_dqdPE7, minv_block_in_R1_C2_dqdPE7, minv_block_in_R2_C2_dqdPE7, minv_block_in_R3_C2_dqdPE7, minv_block_in_R4_C2_dqdPE7, minv_block_in_R5_C2_dqdPE7, minv_block_in_R6_C2_dqdPE7, minv_block_in_R7_C2_dqdPE7, minv_block_in_R1_C3_dqdPE7, minv_block_in_R2_C3_dqdPE7, minv_block_in_R3_C3_dqdPE7, minv_block_in_R4_C3_dqdPE7, minv_block_in_R5_C3_dqdPE7, minv_block_in_R6_C3_dqdPE7, minv_block_in_R7_C3_dqdPE7, minv_block_in_R1_C4_dqdPE7, minv_block_in_R2_C4_dqdPE7, minv_block_in_R3_C4_dqdPE7, minv_block_in_R4_C4_dqdPE7, minv_block_in_R5_C4_dqdPE7, minv_block_in_R6_C4_dqdPE7, minv_block_in_R7_C4_dqdPE7, minv_block_in_R1_C5_dqdPE7, minv_block_in_R2_C5_dqdPE7, minv_block_in_R3_C5_dqdPE7, minv_block_in_R4_C5_dqdPE7, minv_block_in_R5_C5_dqdPE7, minv_block_in_R6_C5_dqdPE7, minv_block_in_R7_C5_dqdPE7, minv_block_in_R1_C6_dqdPE7, minv_block_in_R2_C6_dqdPE7, minv_block_in_R3_C6_dqdPE7, minv_block_in_R4_C6_dqdPE7, minv_block_in_R5_C6_dqdPE7, minv_block_in_R6_C6_dqdPE7, minv_block_in_R7_C6_dqdPE7, minv_block_in_R1_C7_dqdPE7, minv_block_in_R2_C7_dqdPE7, minv_block_in_R3_C7_dqdPE7, minv_block_in_R4_C7_dqdPE7, minv_block_in_R5_C7_dqdPE7, minv_block_in_R6_C7_dqdPE7, minv_block_in_R7_C7_dqdPE7, dtau_vec_in_R1_dqdPE1, dtau_vec_in_R2_dqdPE1, dtau_vec_in_R3_dqdPE1, dtau_vec_in_R4_dqdPE1, dtau_vec_in_R5_dqdPE1, dtau_vec_in_R6_dqdPE1, dtau_vec_in_R7_dqdPE1, dtau_vec_in_R1_dqdPE2, dtau_vec_in_R2_dqdPE2, dtau_vec_in_R3_dqdPE2, dtau_vec_in_R4_dqdPE2, dtau_vec_in_R5_dqdPE2, dtau_vec_in_R6_dqdPE2, dtau_vec_in_R7_dqdPE2, dtau_vec_in_R1_dqdPE3, dtau_vec_in_R2_dqdPE3, dtau_vec_in_R3_dqdPE3, dtau_vec_in_R4_dqdPE3, dtau_vec_in_R5_dqdPE3, dtau_vec_in_R6_dqdPE3, dtau_vec_in_R7_dqdPE3, dtau_vec_in_R1_dqdPE4, dtau_vec_in_R2_dqdPE4, dtau_vec_in_R3_dqdPE4, dtau_vec_in_R4_dqdPE4, dtau_vec_in_R5_dqdPE4, dtau_vec_in_R6_dqdPE4, dtau_vec_in_R7_dqdPE4, dtau_vec_in_R1_dqdPE5, dtau_vec_in_R2_dqdPE5, dtau_vec_in_R3_dqdPE5, dtau_vec_in_R4_dqdPE5, dtau_vec_in_R5_dqdPE5, dtau_vec_in_R6_dqdPE5, dtau_vec_in_R7_dqdPE5, dtau_vec_in_R1_dqdPE6, dtau_vec_in_R2_dqdPE6, dtau_vec_in_R3_dqdPE6, dtau_vec_in_R4_dqdPE6, dtau_vec_in_R5_dqdPE6, dtau_vec_in_R6_dqdPE6, dtau_vec_in_R7_dqdPE6, dtau_vec_in_R1_dqdPE7, dtau_vec_in_R2_dqdPE7, dtau_vec_in_R3_dqdPE7, dtau_vec_in_R4_dqdPE7, dtau_vec_in_R5_dqdPE7, dtau_vec_in_R6_dqdPE7, dtau_vec_in_R7_dqdPE7,
        output_ready, output_ready_minv, tau_curr_out_rnea,
        f_upd_prev_vec_out_AX_rnea, f_upd_prev_vec_out_AY_rnea, f_upd_prev_vec_out_AZ_rnea, f_upd_prev_vec_out_LX_rnea, f_upd_prev_vec_out_LY_rnea, f_upd_prev_vec_out_LZ_rnea,
        dtau_curr_out_dqPE1, dtau_curr_out_dqPE2, dtau_curr_out_dqPE3, dtau_curr_out_dqPE4, dtau_curr_out_dqPE5, dtau_curr_out_dqPE6, dtau_curr_out_dqPE7, dtau_curr_out_dqdPE1, dtau_curr_out_dqdPE2, dtau_curr_out_dqdPE3, dtau_curr_out_dqdPE4, dtau_curr_out_dqdPE5, dtau_curr_out_dqdPE6, dtau_curr_out_dqdPE7, dfdq_upd_prev_vec_out_AX_dqPE1, dfdq_upd_prev_vec_out_AY_dqPE1, dfdq_upd_prev_vec_out_AZ_dqPE1, dfdq_upd_prev_vec_out_LX_dqPE1, dfdq_upd_prev_vec_out_LY_dqPE1, dfdq_upd_prev_vec_out_LZ_dqPE1, dfdq_upd_prev_vec_out_AX_dqPE2, dfdq_upd_prev_vec_out_AY_dqPE2, dfdq_upd_prev_vec_out_AZ_dqPE2, dfdq_upd_prev_vec_out_LX_dqPE2, dfdq_upd_prev_vec_out_LY_dqPE2, dfdq_upd_prev_vec_out_LZ_dqPE2, dfdq_upd_prev_vec_out_AX_dqPE3, dfdq_upd_prev_vec_out_AY_dqPE3, dfdq_upd_prev_vec_out_AZ_dqPE3, dfdq_upd_prev_vec_out_LX_dqPE3, dfdq_upd_prev_vec_out_LY_dqPE3, dfdq_upd_prev_vec_out_LZ_dqPE3, dfdq_upd_prev_vec_out_AX_dqPE4, dfdq_upd_prev_vec_out_AY_dqPE4, dfdq_upd_prev_vec_out_AZ_dqPE4, dfdq_upd_prev_vec_out_LX_dqPE4, dfdq_upd_prev_vec_out_LY_dqPE4, dfdq_upd_prev_vec_out_LZ_dqPE4, dfdq_upd_prev_vec_out_AX_dqPE5, dfdq_upd_prev_vec_out_AY_dqPE5, dfdq_upd_prev_vec_out_AZ_dqPE5, dfdq_upd_prev_vec_out_LX_dqPE5, dfdq_upd_prev_vec_out_LY_dqPE5, dfdq_upd_prev_vec_out_LZ_dqPE5, dfdq_upd_prev_vec_out_AX_dqPE6, dfdq_upd_prev_vec_out_AY_dqPE6, dfdq_upd_prev_vec_out_AZ_dqPE6, dfdq_upd_prev_vec_out_LX_dqPE6, dfdq_upd_prev_vec_out_LY_dqPE6, dfdq_upd_prev_vec_out_LZ_dqPE6, dfdq_upd_prev_vec_out_AX_dqPE7, dfdq_upd_prev_vec_out_AY_dqPE7, dfdq_upd_prev_vec_out_AZ_dqPE7, dfdq_upd_prev_vec_out_LX_dqPE7, dfdq_upd_prev_vec_out_LY_dqPE7, dfdq_upd_prev_vec_out_LZ_dqPE7, dfdqd_upd_prev_vec_out_AX_dqdPE1, dfdqd_upd_prev_vec_out_AY_dqdPE1, dfdqd_upd_prev_vec_out_AZ_dqdPE1, dfdqd_upd_prev_vec_out_LX_dqdPE1, dfdqd_upd_prev_vec_out_LY_dqdPE1, dfdqd_upd_prev_vec_out_LZ_dqdPE1, dfdqd_upd_prev_vec_out_AX_dqdPE2, dfdqd_upd_prev_vec_out_AY_dqdPE2, dfdqd_upd_prev_vec_out_AZ_dqdPE2, dfdqd_upd_prev_vec_out_LX_dqdPE2, dfdqd_upd_prev_vec_out_LY_dqdPE2, dfdqd_upd_prev_vec_out_LZ_dqdPE2, dfdqd_upd_prev_vec_out_AX_dqdPE3, dfdqd_upd_prev_vec_out_AY_dqdPE3, dfdqd_upd_prev_vec_out_AZ_dqdPE3, dfdqd_upd_prev_vec_out_LX_dqdPE3, dfdqd_upd_prev_vec_out_LY_dqdPE3, dfdqd_upd_prev_vec_out_LZ_dqdPE3, dfdqd_upd_prev_vec_out_AX_dqdPE4, dfdqd_upd_prev_vec_out_AY_dqdPE4, dfdqd_upd_prev_vec_out_AZ_dqdPE4, dfdqd_upd_prev_vec_out_LX_dqdPE4, dfdqd_upd_prev_vec_out_LY_dqdPE4, dfdqd_upd_prev_vec_out_LZ_dqdPE4, dfdqd_upd_prev_vec_out_AX_dqdPE5, dfdqd_upd_prev_vec_out_AY_dqdPE5, dfdqd_upd_prev_vec_out_AZ_dqdPE5, dfdqd_upd_prev_vec_out_LX_dqdPE5, dfdqd_upd_prev_vec_out_LY_dqdPE5, dfdqd_upd_prev_vec_out_LZ_dqdPE5, dfdqd_upd_prev_vec_out_AX_dqdPE6, dfdqd_upd_prev_vec_out_AY_dqdPE6, dfdqd_upd_prev_vec_out_AZ_dqdPE6, dfdqd_upd_prev_vec_out_LX_dqdPE6, dfdqd_upd_prev_vec_out_LY_dqdPE6, dfdqd_upd_prev_vec_out_LZ_dqdPE6, dfdqd_upd_prev_vec_out_AX_dqdPE7, dfdqd_upd_prev_vec_out_AY_dqdPE7, dfdqd_upd_prev_vec_out_AZ_dqdPE7, dfdqd_upd_prev_vec_out_LX_dqdPE7, dfdqd_upd_prev_vec_out_LY_dqdPE7, dfdqd_upd_prev_vec_out_LZ_dqdPE7,
        minv_vec_out_R1_dqdPE1, minv_vec_out_R2_dqdPE1, minv_vec_out_R3_dqdPE1, minv_vec_out_R4_dqdPE1, minv_vec_out_R5_dqdPE1, minv_vec_out_R6_dqdPE1, minv_vec_out_R7_dqdPE1, minv_vec_out_R1_dqdPE2, minv_vec_out_R2_dqdPE2, minv_vec_out_R3_dqdPE2, minv_vec_out_R4_dqdPE2, minv_vec_out_R5_dqdPE2, minv_vec_out_R6_dqdPE2, minv_vec_out_R7_dqdPE2, minv_vec_out_R1_dqdPE3, minv_vec_out_R2_dqdPE3, minv_vec_out_R3_dqdPE3, minv_vec_out_R4_dqdPE3, minv_vec_out_R5_dqdPE3, minv_vec_out_R6_dqdPE3, minv_vec_out_R7_dqdPE3, minv_vec_out_R1_dqdPE4, minv_vec_out_R2_dqdPE4, minv_vec_out_R3_dqdPE4, minv_vec_out_R4_dqdPE4, minv_vec_out_R5_dqdPE4, minv_vec_out_R6_dqdPE4, minv_vec_out_R7_dqdPE4, minv_vec_out_R1_dqdPE5, minv_vec_out_R2_dqdPE5, minv_vec_out_R3_dqdPE5, minv_vec_out_R4_dqdPE5, minv_vec_out_R5_dqdPE5, minv_vec_out_R6_dqdPE5, minv_vec_out_R7_dqdPE5, minv_vec_out_R1_dqdPE6, minv_vec_out_R2_dqdPE6, minv_vec_out_R3_dqdPE6, minv_vec_out_R4_dqdPE6, minv_vec_out_R5_dqdPE6, minv_vec_out_R6_dqdPE6, minv_vec_out_R7_dqdPE6, minv_vec_out_R1_dqdPE7, minv_vec_out_R2_dqdPE7, minv_vec_out_R3_dqdPE7, minv_vec_out_R4_dqdPE7, minv_vec_out_R5_dqdPE7, minv_vec_out_R6_dqdPE7, minv_vec_out_R7_dqdPE7
    ) CF (
        get_data, get_data_minv, link_in_rnea, sinq_val_in_rnea, cosq_val_in_rnea,
        f_upd_curr_vec_in_AX_rnea, f_upd_curr_vec_in_AY_rnea, f_upd_curr_vec_in_AZ_rnea, f_upd_curr_vec_in_LX_rnea, f_upd_curr_vec_in_LY_rnea, f_upd_curr_vec_in_LZ_rnea, f_prev_vec_in_AX_rnea, f_prev_vec_in_AY_rnea, f_prev_vec_in_AZ_rnea, f_prev_vec_in_LX_rnea, f_prev_vec_in_LY_rnea, f_prev_vec_in_LZ_rnea,
        link_in_dqPE1, link_in_dqPE2, link_in_dqPE3, link_in_dqPE4, link_in_dqPE5, link_in_dqPE6, link_in_dqPE7, link_in_dqdPE1, link_in_dqdPE2, link_in_dqdPE3, link_in_dqdPE4, link_in_dqdPE5, link_in_dqdPE6, link_in_dqdPE7, derv_in_dqPE1, derv_in_dqPE2, derv_in_dqPE3, derv_in_dqPE4, derv_in_dqPE5, derv_in_dqPE6, derv_in_dqPE7, derv_in_dqdPE1, derv_in_dqdPE2, derv_in_dqdPE3, derv_in_dqdPE4, derv_in_dqdPE5, derv_in_dqdPE6, derv_in_dqdPE7,
        sinq_val_in_dqPE1, sinq_val_in_dqPE2, sinq_val_in_dqPE3, sinq_val_in_dqPE4, sinq_val_in_dqPE5, sinq_val_in_dqPE6, sinq_val_in_dqPE7, sinq_val_in_dqdPE1, sinq_val_in_dqdPE2, sinq_val_in_dqdPE3, sinq_val_in_dqdPE4, sinq_val_in_dqdPE5, sinq_val_in_dqdPE6, sinq_val_in_dqdPE7, cosq_val_in_dqPE1, cosq_val_in_dqPE2, cosq_val_in_dqPE3, cosq_val_in_dqPE4, cosq_val_in_dqPE5, cosq_val_in_dqPE6, cosq_val_in_dqPE7, cosq_val_in_dqdPE1, cosq_val_in_dqdPE2, cosq_val_in_dqdPE3, cosq_val_in_dqdPE4, cosq_val_in_dqdPE5, cosq_val_in_dqdPE6, cosq_val_in_dqdPE7,
        f_upd_curr_vec_in_AX_dqPE1, f_upd_curr_vec_in_AY_dqPE1, f_upd_curr_vec_in_AZ_dqPE1, f_upd_curr_vec_in_LX_dqPE1, f_upd_curr_vec_in_LY_dqPE1, f_upd_curr_vec_in_LZ_dqPE1, f_upd_curr_vec_in_AX_dqPE2, f_upd_curr_vec_in_AY_dqPE2, f_upd_curr_vec_in_AZ_dqPE2, f_upd_curr_vec_in_LX_dqPE2, f_upd_curr_vec_in_LY_dqPE2, f_upd_curr_vec_in_LZ_dqPE2, f_upd_curr_vec_in_AX_dqPE3, f_upd_curr_vec_in_AY_dqPE3, f_upd_curr_vec_in_AZ_dqPE3, f_upd_curr_vec_in_LX_dqPE3, f_upd_curr_vec_in_LY_dqPE3, f_upd_curr_vec_in_LZ_dqPE3, f_upd_curr_vec_in_AX_dqPE4, f_upd_curr_vec_in_AY_dqPE4, f_upd_curr_vec_in_AZ_dqPE4, f_upd_curr_vec_in_LX_dqPE4, f_upd_curr_vec_in_LY_dqPE4, f_upd_curr_vec_in_LZ_dqPE4, f_upd_curr_vec_in_AX_dqPE5, f_upd_curr_vec_in_AY_dqPE5, f_upd_curr_vec_in_AZ_dqPE5, f_upd_curr_vec_in_LX_dqPE5, f_upd_curr_vec_in_LY_dqPE5, f_upd_curr_vec_in_LZ_dqPE5, f_upd_curr_vec_in_AX_dqPE6, f_upd_curr_vec_in_AY_dqPE6, f_upd_curr_vec_in_AZ_dqPE6, f_upd_curr_vec_in_LX_dqPE6, f_upd_curr_vec_in_LY_dqPE6, f_upd_curr_vec_in_LZ_dqPE6, f_upd_curr_vec_in_AX_dqPE7, f_upd_curr_vec_in_AY_dqPE7, f_upd_curr_vec_in_AZ_dqPE7, f_upd_curr_vec_in_LX_dqPE7, f_upd_curr_vec_in_LY_dqPE7, f_upd_curr_vec_in_LZ_dqPE7, dfdq_prev_vec_in_AX_dqPE1, dfdq_prev_vec_in_AY_dqPE1, dfdq_prev_vec_in_AZ_dqPE1, dfdq_prev_vec_in_LX_dqPE1, dfdq_prev_vec_in_LY_dqPE1, dfdq_prev_vec_in_LZ_dqPE1, dfdq_prev_vec_in_AX_dqPE2, dfdq_prev_vec_in_AY_dqPE2, dfdq_prev_vec_in_AZ_dqPE2, dfdq_prev_vec_in_LX_dqPE2, dfdq_prev_vec_in_LY_dqPE2, dfdq_prev_vec_in_LZ_dqPE2, dfdq_prev_vec_in_AX_dqPE3, dfdq_prev_vec_in_AY_dqPE3, dfdq_prev_vec_in_AZ_dqPE3, dfdq_prev_vec_in_LX_dqPE3, dfdq_prev_vec_in_LY_dqPE3, dfdq_prev_vec_in_LZ_dqPE3, dfdq_prev_vec_in_AX_dqPE4, dfdq_prev_vec_in_AY_dqPE4, dfdq_prev_vec_in_AZ_dqPE4, dfdq_prev_vec_in_LX_dqPE4, dfdq_prev_vec_in_LY_dqPE4, dfdq_prev_vec_in_LZ_dqPE4, dfdq_prev_vec_in_AX_dqPE5, dfdq_prev_vec_in_AY_dqPE5, dfdq_prev_vec_in_AZ_dqPE5, dfdq_prev_vec_in_LX_dqPE5, dfdq_prev_vec_in_LY_dqPE5, dfdq_prev_vec_in_LZ_dqPE5, dfdq_prev_vec_in_AX_dqPE6, dfdq_prev_vec_in_AY_dqPE6, dfdq_prev_vec_in_AZ_dqPE6, dfdq_prev_vec_in_LX_dqPE6, dfdq_prev_vec_in_LY_dqPE6, dfdq_prev_vec_in_LZ_dqPE6, dfdq_prev_vec_in_AX_dqPE7, dfdq_prev_vec_in_AY_dqPE7, dfdq_prev_vec_in_AZ_dqPE7, dfdq_prev_vec_in_LX_dqPE7, dfdq_prev_vec_in_LY_dqPE7, dfdq_prev_vec_in_LZ_dqPE7, dfdq_upd_curr_vec_in_AX_dqPE1, dfdq_upd_curr_vec_in_AY_dqPE1, dfdq_upd_curr_vec_in_AZ_dqPE1, dfdq_upd_curr_vec_in_LX_dqPE1, dfdq_upd_curr_vec_in_LY_dqPE1, dfdq_upd_curr_vec_in_LZ_dqPE1, dfdq_upd_curr_vec_in_AX_dqPE2, dfdq_upd_curr_vec_in_AY_dqPE2, dfdq_upd_curr_vec_in_AZ_dqPE2, dfdq_upd_curr_vec_in_LX_dqPE2, dfdq_upd_curr_vec_in_LY_dqPE2, dfdq_upd_curr_vec_in_LZ_dqPE2, dfdq_upd_curr_vec_in_AX_dqPE3, dfdq_upd_curr_vec_in_AY_dqPE3, dfdq_upd_curr_vec_in_AZ_dqPE3, dfdq_upd_curr_vec_in_LX_dqPE3, dfdq_upd_curr_vec_in_LY_dqPE3, dfdq_upd_curr_vec_in_LZ_dqPE3, dfdq_upd_curr_vec_in_AX_dqPE4, dfdq_upd_curr_vec_in_AY_dqPE4, dfdq_upd_curr_vec_in_AZ_dqPE4, dfdq_upd_curr_vec_in_LX_dqPE4, dfdq_upd_curr_vec_in_LY_dqPE4, dfdq_upd_curr_vec_in_LZ_dqPE4, dfdq_upd_curr_vec_in_AX_dqPE5, dfdq_upd_curr_vec_in_AY_dqPE5, dfdq_upd_curr_vec_in_AZ_dqPE5, dfdq_upd_curr_vec_in_LX_dqPE5, dfdq_upd_curr_vec_in_LY_dqPE5, dfdq_upd_curr_vec_in_LZ_dqPE5, dfdq_upd_curr_vec_in_AX_dqPE6, dfdq_upd_curr_vec_in_AY_dqPE6, dfdq_upd_curr_vec_in_AZ_dqPE6, dfdq_upd_curr_vec_in_LX_dqPE6, dfdq_upd_curr_vec_in_LY_dqPE6, dfdq_upd_curr_vec_in_LZ_dqPE6, dfdq_upd_curr_vec_in_AX_dqPE7, dfdq_upd_curr_vec_in_AY_dqPE7, dfdq_upd_curr_vec_in_AZ_dqPE7, dfdq_upd_curr_vec_in_LX_dqPE7, dfdq_upd_curr_vec_in_LY_dqPE7, dfdq_upd_curr_vec_in_LZ_dqPE7, dfdqd_prev_vec_in_AX_dqdPE1, dfdqd_prev_vec_in_AY_dqdPE1, dfdqd_prev_vec_in_AZ_dqdPE1, dfdqd_prev_vec_in_LX_dqdPE1, dfdqd_prev_vec_in_LY_dqdPE1, dfdqd_prev_vec_in_LZ_dqdPE1, dfdqd_prev_vec_in_AX_dqdPE2, dfdqd_prev_vec_in_AY_dqdPE2, dfdqd_prev_vec_in_AZ_dqdPE2, dfdqd_prev_vec_in_LX_dqdPE2, dfdqd_prev_vec_in_LY_dqdPE2, dfdqd_prev_vec_in_LZ_dqdPE2, dfdqd_prev_vec_in_AX_dqdPE3, dfdqd_prev_vec_in_AY_dqdPE3, dfdqd_prev_vec_in_AZ_dqdPE3, dfdqd_prev_vec_in_LX_dqdPE3, dfdqd_prev_vec_in_LY_dqdPE3, dfdqd_prev_vec_in_LZ_dqdPE3, dfdqd_prev_vec_in_AX_dqdPE4, dfdqd_prev_vec_in_AY_dqdPE4, dfdqd_prev_vec_in_AZ_dqdPE4, dfdqd_prev_vec_in_LX_dqdPE4, dfdqd_prev_vec_in_LY_dqdPE4, dfdqd_prev_vec_in_LZ_dqdPE4, dfdqd_prev_vec_in_AX_dqdPE5, dfdqd_prev_vec_in_AY_dqdPE5, dfdqd_prev_vec_in_AZ_dqdPE5, dfdqd_prev_vec_in_LX_dqdPE5, dfdqd_prev_vec_in_LY_dqdPE5, dfdqd_prev_vec_in_LZ_dqdPE5, dfdqd_prev_vec_in_AX_dqdPE6, dfdqd_prev_vec_in_AY_dqdPE6, dfdqd_prev_vec_in_AZ_dqdPE6, dfdqd_prev_vec_in_LX_dqdPE6, dfdqd_prev_vec_in_LY_dqdPE6, dfdqd_prev_vec_in_LZ_dqdPE6, dfdqd_prev_vec_in_AX_dqdPE7, dfdqd_prev_vec_in_AY_dqdPE7, dfdqd_prev_vec_in_AZ_dqdPE7, dfdqd_prev_vec_in_LX_dqdPE7, dfdqd_prev_vec_in_LY_dqdPE7, dfdqd_prev_vec_in_LZ_dqdPE7, dfdqd_upd_curr_vec_in_AX_dqdPE1, dfdqd_upd_curr_vec_in_AY_dqdPE1, dfdqd_upd_curr_vec_in_AZ_dqdPE1, dfdqd_upd_curr_vec_in_LX_dqdPE1, dfdqd_upd_curr_vec_in_LY_dqdPE1, dfdqd_upd_curr_vec_in_LZ_dqdPE1, dfdqd_upd_curr_vec_in_AX_dqdPE2, dfdqd_upd_curr_vec_in_AY_dqdPE2, dfdqd_upd_curr_vec_in_AZ_dqdPE2, dfdqd_upd_curr_vec_in_LX_dqdPE2, dfdqd_upd_curr_vec_in_LY_dqdPE2, dfdqd_upd_curr_vec_in_LZ_dqdPE2, dfdqd_upd_curr_vec_in_AX_dqdPE3, dfdqd_upd_curr_vec_in_AY_dqdPE3, dfdqd_upd_curr_vec_in_AZ_dqdPE3, dfdqd_upd_curr_vec_in_LX_dqdPE3, dfdqd_upd_curr_vec_in_LY_dqdPE3, dfdqd_upd_curr_vec_in_LZ_dqdPE3, dfdqd_upd_curr_vec_in_AX_dqdPE4, dfdqd_upd_curr_vec_in_AY_dqdPE4, dfdqd_upd_curr_vec_in_AZ_dqdPE4, dfdqd_upd_curr_vec_in_LX_dqdPE4, dfdqd_upd_curr_vec_in_LY_dqdPE4, dfdqd_upd_curr_vec_in_LZ_dqdPE4, dfdqd_upd_curr_vec_in_AX_dqdPE5, dfdqd_upd_curr_vec_in_AY_dqdPE5, dfdqd_upd_curr_vec_in_AZ_dqdPE5, dfdqd_upd_curr_vec_in_LX_dqdPE5, dfdqd_upd_curr_vec_in_LY_dqdPE5, dfdqd_upd_curr_vec_in_LZ_dqdPE5, dfdqd_upd_curr_vec_in_AX_dqdPE6, dfdqd_upd_curr_vec_in_AY_dqdPE6, dfdqd_upd_curr_vec_in_AZ_dqdPE6, dfdqd_upd_curr_vec_in_LX_dqdPE6, dfdqd_upd_curr_vec_in_LY_dqdPE6, dfdqd_upd_curr_vec_in_LZ_dqdPE6, dfdqd_upd_curr_vec_in_AX_dqdPE7, dfdqd_upd_curr_vec_in_AY_dqdPE7, dfdqd_upd_curr_vec_in_AZ_dqdPE7, dfdqd_upd_curr_vec_in_LX_dqdPE7, dfdqd_upd_curr_vec_in_LY_dqdPE7, dfdqd_upd_curr_vec_in_LZ_dqdPE7,
        minv_block_in_R1_C1_dqdPE1, minv_block_in_R2_C1_dqdPE1, minv_block_in_R3_C1_dqdPE1, minv_block_in_R4_C1_dqdPE1, minv_block_in_R5_C1_dqdPE1, minv_block_in_R6_C1_dqdPE1, minv_block_in_R7_C1_dqdPE1, minv_block_in_R1_C2_dqdPE1, minv_block_in_R2_C2_dqdPE1, minv_block_in_R3_C2_dqdPE1, minv_block_in_R4_C2_dqdPE1, minv_block_in_R5_C2_dqdPE1, minv_block_in_R6_C2_dqdPE1, minv_block_in_R7_C2_dqdPE1, minv_block_in_R1_C3_dqdPE1, minv_block_in_R2_C3_dqdPE1, minv_block_in_R3_C3_dqdPE1, minv_block_in_R4_C3_dqdPE1, minv_block_in_R5_C3_dqdPE1, minv_block_in_R6_C3_dqdPE1, minv_block_in_R7_C3_dqdPE1, minv_block_in_R1_C4_dqdPE1, minv_block_in_R2_C4_dqdPE1, minv_block_in_R3_C4_dqdPE1, minv_block_in_R4_C4_dqdPE1, minv_block_in_R5_C4_dqdPE1, minv_block_in_R6_C4_dqdPE1, minv_block_in_R7_C4_dqdPE1, minv_block_in_R1_C5_dqdPE1, minv_block_in_R2_C5_dqdPE1, minv_block_in_R3_C5_dqdPE1, minv_block_in_R4_C5_dqdPE1, minv_block_in_R5_C5_dqdPE1, minv_block_in_R6_C5_dqdPE1, minv_block_in_R7_C5_dqdPE1, minv_block_in_R1_C6_dqdPE1, minv_block_in_R2_C6_dqdPE1, minv_block_in_R3_C6_dqdPE1, minv_block_in_R4_C6_dqdPE1, minv_block_in_R5_C6_dqdPE1, minv_block_in_R6_C6_dqdPE1, minv_block_in_R7_C6_dqdPE1, minv_block_in_R1_C7_dqdPE1, minv_block_in_R2_C7_dqdPE1, minv_block_in_R3_C7_dqdPE1, minv_block_in_R4_C7_dqdPE1, minv_block_in_R5_C7_dqdPE1, minv_block_in_R6_C7_dqdPE1, minv_block_in_R7_C7_dqdPE1, minv_block_in_R1_C1_dqdPE2, minv_block_in_R2_C1_dqdPE2, minv_block_in_R3_C1_dqdPE2, minv_block_in_R4_C1_dqdPE2, minv_block_in_R5_C1_dqdPE2, minv_block_in_R6_C1_dqdPE2, minv_block_in_R7_C1_dqdPE2, minv_block_in_R1_C2_dqdPE2, minv_block_in_R2_C2_dqdPE2, minv_block_in_R3_C2_dqdPE2, minv_block_in_R4_C2_dqdPE2, minv_block_in_R5_C2_dqdPE2, minv_block_in_R6_C2_dqdPE2, minv_block_in_R7_C2_dqdPE2, minv_block_in_R1_C3_dqdPE2, minv_block_in_R2_C3_dqdPE2, minv_block_in_R3_C3_dqdPE2, minv_block_in_R4_C3_dqdPE2, minv_block_in_R5_C3_dqdPE2, minv_block_in_R6_C3_dqdPE2, minv_block_in_R7_C3_dqdPE2, minv_block_in_R1_C4_dqdPE2, minv_block_in_R2_C4_dqdPE2, minv_block_in_R3_C4_dqdPE2, minv_block_in_R4_C4_dqdPE2, minv_block_in_R5_C4_dqdPE2, minv_block_in_R6_C4_dqdPE2, minv_block_in_R7_C4_dqdPE2, minv_block_in_R1_C5_dqdPE2, minv_block_in_R2_C5_dqdPE2, minv_block_in_R3_C5_dqdPE2, minv_block_in_R4_C5_dqdPE2, minv_block_in_R5_C5_dqdPE2, minv_block_in_R6_C5_dqdPE2, minv_block_in_R7_C5_dqdPE2, minv_block_in_R1_C6_dqdPE2, minv_block_in_R2_C6_dqdPE2, minv_block_in_R3_C6_dqdPE2, minv_block_in_R4_C6_dqdPE2, minv_block_in_R5_C6_dqdPE2, minv_block_in_R6_C6_dqdPE2, minv_block_in_R7_C6_dqdPE2, minv_block_in_R1_C7_dqdPE2, minv_block_in_R2_C7_dqdPE2, minv_block_in_R3_C7_dqdPE2, minv_block_in_R4_C7_dqdPE2, minv_block_in_R5_C7_dqdPE2, minv_block_in_R6_C7_dqdPE2, minv_block_in_R7_C7_dqdPE2, minv_block_in_R1_C1_dqdPE3, minv_block_in_R2_C1_dqdPE3, minv_block_in_R3_C1_dqdPE3, minv_block_in_R4_C1_dqdPE3, minv_block_in_R5_C1_dqdPE3, minv_block_in_R6_C1_dqdPE3, minv_block_in_R7_C1_dqdPE3, minv_block_in_R1_C2_dqdPE3, minv_block_in_R2_C2_dqdPE3, minv_block_in_R3_C2_dqdPE3, minv_block_in_R4_C2_dqdPE3, minv_block_in_R5_C2_dqdPE3, minv_block_in_R6_C2_dqdPE3, minv_block_in_R7_C2_dqdPE3, minv_block_in_R1_C3_dqdPE3, minv_block_in_R2_C3_dqdPE3, minv_block_in_R3_C3_dqdPE3, minv_block_in_R4_C3_dqdPE3, minv_block_in_R5_C3_dqdPE3, minv_block_in_R6_C3_dqdPE3, minv_block_in_R7_C3_dqdPE3, minv_block_in_R1_C4_dqdPE3, minv_block_in_R2_C4_dqdPE3, minv_block_in_R3_C4_dqdPE3, minv_block_in_R4_C4_dqdPE3, minv_block_in_R5_C4_dqdPE3, minv_block_in_R6_C4_dqdPE3, minv_block_in_R7_C4_dqdPE3, minv_block_in_R1_C5_dqdPE3, minv_block_in_R2_C5_dqdPE3, minv_block_in_R3_C5_dqdPE3, minv_block_in_R4_C5_dqdPE3, minv_block_in_R5_C5_dqdPE3, minv_block_in_R6_C5_dqdPE3, minv_block_in_R7_C5_dqdPE3, minv_block_in_R1_C6_dqdPE3, minv_block_in_R2_C6_dqdPE3, minv_block_in_R3_C6_dqdPE3, minv_block_in_R4_C6_dqdPE3, minv_block_in_R5_C6_dqdPE3, minv_block_in_R6_C6_dqdPE3, minv_block_in_R7_C6_dqdPE3, minv_block_in_R1_C7_dqdPE3, minv_block_in_R2_C7_dqdPE3, minv_block_in_R3_C7_dqdPE3, minv_block_in_R4_C7_dqdPE3, minv_block_in_R5_C7_dqdPE3, minv_block_in_R6_C7_dqdPE3, minv_block_in_R7_C7_dqdPE3, minv_block_in_R1_C1_dqdPE4, minv_block_in_R2_C1_dqdPE4, minv_block_in_R3_C1_dqdPE4, minv_block_in_R4_C1_dqdPE4, minv_block_in_R5_C1_dqdPE4, minv_block_in_R6_C1_dqdPE4, minv_block_in_R7_C1_dqdPE4, minv_block_in_R1_C2_dqdPE4, minv_block_in_R2_C2_dqdPE4, minv_block_in_R3_C2_dqdPE4, minv_block_in_R4_C2_dqdPE4, minv_block_in_R5_C2_dqdPE4, minv_block_in_R6_C2_dqdPE4, minv_block_in_R7_C2_dqdPE4, minv_block_in_R1_C3_dqdPE4, minv_block_in_R2_C3_dqdPE4, minv_block_in_R3_C3_dqdPE4, minv_block_in_R4_C3_dqdPE4, minv_block_in_R5_C3_dqdPE4, minv_block_in_R6_C3_dqdPE4, minv_block_in_R7_C3_dqdPE4, minv_block_in_R1_C4_dqdPE4, minv_block_in_R2_C4_dqdPE4, minv_block_in_R3_C4_dqdPE4, minv_block_in_R4_C4_dqdPE4, minv_block_in_R5_C4_dqdPE4, minv_block_in_R6_C4_dqdPE4, minv_block_in_R7_C4_dqdPE4, minv_block_in_R1_C5_dqdPE4, minv_block_in_R2_C5_dqdPE4, minv_block_in_R3_C5_dqdPE4, minv_block_in_R4_C5_dqdPE4, minv_block_in_R5_C5_dqdPE4, minv_block_in_R6_C5_dqdPE4, minv_block_in_R7_C5_dqdPE4, minv_block_in_R1_C6_dqdPE4, minv_block_in_R2_C6_dqdPE4, minv_block_in_R3_C6_dqdPE4, minv_block_in_R4_C6_dqdPE4, minv_block_in_R5_C6_dqdPE4, minv_block_in_R6_C6_dqdPE4, minv_block_in_R7_C6_dqdPE4, minv_block_in_R1_C7_dqdPE4, minv_block_in_R2_C7_dqdPE4, minv_block_in_R3_C7_dqdPE4, minv_block_in_R4_C7_dqdPE4, minv_block_in_R5_C7_dqdPE4, minv_block_in_R6_C7_dqdPE4, minv_block_in_R7_C7_dqdPE4, minv_block_in_R1_C1_dqdPE5, minv_block_in_R2_C1_dqdPE5, minv_block_in_R3_C1_dqdPE5, minv_block_in_R4_C1_dqdPE5, minv_block_in_R5_C1_dqdPE5, minv_block_in_R6_C1_dqdPE5, minv_block_in_R7_C1_dqdPE5, minv_block_in_R1_C2_dqdPE5, minv_block_in_R2_C2_dqdPE5, minv_block_in_R3_C2_dqdPE5, minv_block_in_R4_C2_dqdPE5, minv_block_in_R5_C2_dqdPE5, minv_block_in_R6_C2_dqdPE5, minv_block_in_R7_C2_dqdPE5, minv_block_in_R1_C3_dqdPE5, minv_block_in_R2_C3_dqdPE5, minv_block_in_R3_C3_dqdPE5, minv_block_in_R4_C3_dqdPE5, minv_block_in_R5_C3_dqdPE5, minv_block_in_R6_C3_dqdPE5, minv_block_in_R7_C3_dqdPE5, minv_block_in_R1_C4_dqdPE5, minv_block_in_R2_C4_dqdPE5, minv_block_in_R3_C4_dqdPE5, minv_block_in_R4_C4_dqdPE5, minv_block_in_R5_C4_dqdPE5, minv_block_in_R6_C4_dqdPE5, minv_block_in_R7_C4_dqdPE5, minv_block_in_R1_C5_dqdPE5, minv_block_in_R2_C5_dqdPE5, minv_block_in_R3_C5_dqdPE5, minv_block_in_R4_C5_dqdPE5, minv_block_in_R5_C5_dqdPE5, minv_block_in_R6_C5_dqdPE5, minv_block_in_R7_C5_dqdPE5, minv_block_in_R1_C6_dqdPE5, minv_block_in_R2_C6_dqdPE5, minv_block_in_R3_C6_dqdPE5, minv_block_in_R4_C6_dqdPE5, minv_block_in_R5_C6_dqdPE5, minv_block_in_R6_C6_dqdPE5, minv_block_in_R7_C6_dqdPE5, minv_block_in_R1_C7_dqdPE5, minv_block_in_R2_C7_dqdPE5, minv_block_in_R3_C7_dqdPE5, minv_block_in_R4_C7_dqdPE5, minv_block_in_R5_C7_dqdPE5, minv_block_in_R6_C7_dqdPE5, minv_block_in_R7_C7_dqdPE5, minv_block_in_R1_C1_dqdPE6, minv_block_in_R2_C1_dqdPE6, minv_block_in_R3_C1_dqdPE6, minv_block_in_R4_C1_dqdPE6, minv_block_in_R5_C1_dqdPE6, minv_block_in_R6_C1_dqdPE6, minv_block_in_R7_C1_dqdPE6, minv_block_in_R1_C2_dqdPE6, minv_block_in_R2_C2_dqdPE6, minv_block_in_R3_C2_dqdPE6, minv_block_in_R4_C2_dqdPE6, minv_block_in_R5_C2_dqdPE6, minv_block_in_R6_C2_dqdPE6, minv_block_in_R7_C2_dqdPE6, minv_block_in_R1_C3_dqdPE6, minv_block_in_R2_C3_dqdPE6, minv_block_in_R3_C3_dqdPE6, minv_block_in_R4_C3_dqdPE6, minv_block_in_R5_C3_dqdPE6, minv_block_in_R6_C3_dqdPE6, minv_block_in_R7_C3_dqdPE6, minv_block_in_R1_C4_dqdPE6, minv_block_in_R2_C4_dqdPE6, minv_block_in_R3_C4_dqdPE6, minv_block_in_R4_C4_dqdPE6, minv_block_in_R5_C4_dqdPE6, minv_block_in_R6_C4_dqdPE6, minv_block_in_R7_C4_dqdPE6, minv_block_in_R1_C5_dqdPE6, minv_block_in_R2_C5_dqdPE6, minv_block_in_R3_C5_dqdPE6, minv_block_in_R4_C5_dqdPE6, minv_block_in_R5_C5_dqdPE6, minv_block_in_R6_C5_dqdPE6, minv_block_in_R7_C5_dqdPE6, minv_block_in_R1_C6_dqdPE6, minv_block_in_R2_C6_dqdPE6, minv_block_in_R3_C6_dqdPE6, minv_block_in_R4_C6_dqdPE6, minv_block_in_R5_C6_dqdPE6, minv_block_in_R6_C6_dqdPE6, minv_block_in_R7_C6_dqdPE6, minv_block_in_R1_C7_dqdPE6, minv_block_in_R2_C7_dqdPE6, minv_block_in_R3_C7_dqdPE6, minv_block_in_R4_C7_dqdPE6, minv_block_in_R5_C7_dqdPE6, minv_block_in_R6_C7_dqdPE6, minv_block_in_R7_C7_dqdPE6, minv_block_in_R1_C1_dqdPE7, minv_block_in_R2_C1_dqdPE7, minv_block_in_R3_C1_dqdPE7, minv_block_in_R4_C1_dqdPE7, minv_block_in_R5_C1_dqdPE7, minv_block_in_R6_C1_dqdPE7, minv_block_in_R7_C1_dqdPE7, minv_block_in_R1_C2_dqdPE7, minv_block_in_R2_C2_dqdPE7, minv_block_in_R3_C2_dqdPE7, minv_block_in_R4_C2_dqdPE7, minv_block_in_R5_C2_dqdPE7, minv_block_in_R6_C2_dqdPE7, minv_block_in_R7_C2_dqdPE7, minv_block_in_R1_C3_dqdPE7, minv_block_in_R2_C3_dqdPE7, minv_block_in_R3_C3_dqdPE7, minv_block_in_R4_C3_dqdPE7, minv_block_in_R5_C3_dqdPE7, minv_block_in_R6_C3_dqdPE7, minv_block_in_R7_C3_dqdPE7, minv_block_in_R1_C4_dqdPE7, minv_block_in_R2_C4_dqdPE7, minv_block_in_R3_C4_dqdPE7, minv_block_in_R4_C4_dqdPE7, minv_block_in_R5_C4_dqdPE7, minv_block_in_R6_C4_dqdPE7, minv_block_in_R7_C4_dqdPE7, minv_block_in_R1_C5_dqdPE7, minv_block_in_R2_C5_dqdPE7, minv_block_in_R3_C5_dqdPE7, minv_block_in_R4_C5_dqdPE7, minv_block_in_R5_C5_dqdPE7, minv_block_in_R6_C5_dqdPE7, minv_block_in_R7_C5_dqdPE7, minv_block_in_R1_C6_dqdPE7, minv_block_in_R2_C6_dqdPE7, minv_block_in_R3_C6_dqdPE7, minv_block_in_R4_C6_dqdPE7, minv_block_in_R5_C6_dqdPE7, minv_block_in_R6_C6_dqdPE7, minv_block_in_R7_C6_dqdPE7, minv_block_in_R1_C7_dqdPE7, minv_block_in_R2_C7_dqdPE7, minv_block_in_R3_C7_dqdPE7, minv_block_in_R4_C7_dqdPE7, minv_block_in_R5_C7_dqdPE7, minv_block_in_R6_C7_dqdPE7, minv_block_in_R7_C7_dqdPE7, dtau_vec_in_R1_dqdPE1, dtau_vec_in_R2_dqdPE1, dtau_vec_in_R3_dqdPE1, dtau_vec_in_R4_dqdPE1, dtau_vec_in_R5_dqdPE1, dtau_vec_in_R6_dqdPE1, dtau_vec_in_R7_dqdPE1, dtau_vec_in_R1_dqdPE2, dtau_vec_in_R2_dqdPE2, dtau_vec_in_R3_dqdPE2, dtau_vec_in_R4_dqdPE2, dtau_vec_in_R5_dqdPE2, dtau_vec_in_R6_dqdPE2, dtau_vec_in_R7_dqdPE2, dtau_vec_in_R1_dqdPE3, dtau_vec_in_R2_dqdPE3, dtau_vec_in_R3_dqdPE3, dtau_vec_in_R4_dqdPE3, dtau_vec_in_R5_dqdPE3, dtau_vec_in_R6_dqdPE3, dtau_vec_in_R7_dqdPE3, dtau_vec_in_R1_dqdPE4, dtau_vec_in_R2_dqdPE4, dtau_vec_in_R3_dqdPE4, dtau_vec_in_R4_dqdPE4, dtau_vec_in_R5_dqdPE4, dtau_vec_in_R6_dqdPE4, dtau_vec_in_R7_dqdPE4, dtau_vec_in_R1_dqdPE5, dtau_vec_in_R2_dqdPE5, dtau_vec_in_R3_dqdPE5, dtau_vec_in_R4_dqdPE5, dtau_vec_in_R5_dqdPE5, dtau_vec_in_R6_dqdPE5, dtau_vec_in_R7_dqdPE5, dtau_vec_in_R1_dqdPE6, dtau_vec_in_R2_dqdPE6, dtau_vec_in_R3_dqdPE6, dtau_vec_in_R4_dqdPE6, dtau_vec_in_R5_dqdPE6, dtau_vec_in_R6_dqdPE6, dtau_vec_in_R7_dqdPE6, dtau_vec_in_R1_dqdPE7, dtau_vec_in_R2_dqdPE7, dtau_vec_in_R3_dqdPE7, dtau_vec_in_R4_dqdPE7, dtau_vec_in_R5_dqdPE7, dtau_vec_in_R6_dqdPE7, dtau_vec_in_R7_dqdPE7,
        output_ready, output_ready_minv, tau_curr_out_rnea,
        f_upd_prev_vec_out_AX_rnea, f_upd_prev_vec_out_AY_rnea, f_upd_prev_vec_out_AZ_rnea, f_upd_prev_vec_out_LX_rnea, f_upd_prev_vec_out_LY_rnea, f_upd_prev_vec_out_LZ_rnea,
        dtau_curr_out_dqPE1, dtau_curr_out_dqPE2, dtau_curr_out_dqPE3, dtau_curr_out_dqPE4, dtau_curr_out_dqPE5, dtau_curr_out_dqPE6, dtau_curr_out_dqPE7, dtau_curr_out_dqdPE1, dtau_curr_out_dqdPE2, dtau_curr_out_dqdPE3, dtau_curr_out_dqdPE4, dtau_curr_out_dqdPE5, dtau_curr_out_dqdPE6, dtau_curr_out_dqdPE7, dfdq_upd_prev_vec_out_AX_dqPE1, dfdq_upd_prev_vec_out_AY_dqPE1, dfdq_upd_prev_vec_out_AZ_dqPE1, dfdq_upd_prev_vec_out_LX_dqPE1, dfdq_upd_prev_vec_out_LY_dqPE1, dfdq_upd_prev_vec_out_LZ_dqPE1, dfdq_upd_prev_vec_out_AX_dqPE2, dfdq_upd_prev_vec_out_AY_dqPE2, dfdq_upd_prev_vec_out_AZ_dqPE2, dfdq_upd_prev_vec_out_LX_dqPE2, dfdq_upd_prev_vec_out_LY_dqPE2, dfdq_upd_prev_vec_out_LZ_dqPE2, dfdq_upd_prev_vec_out_AX_dqPE3, dfdq_upd_prev_vec_out_AY_dqPE3, dfdq_upd_prev_vec_out_AZ_dqPE3, dfdq_upd_prev_vec_out_LX_dqPE3, dfdq_upd_prev_vec_out_LY_dqPE3, dfdq_upd_prev_vec_out_LZ_dqPE3, dfdq_upd_prev_vec_out_AX_dqPE4, dfdq_upd_prev_vec_out_AY_dqPE4, dfdq_upd_prev_vec_out_AZ_dqPE4, dfdq_upd_prev_vec_out_LX_dqPE4, dfdq_upd_prev_vec_out_LY_dqPE4, dfdq_upd_prev_vec_out_LZ_dqPE4, dfdq_upd_prev_vec_out_AX_dqPE5, dfdq_upd_prev_vec_out_AY_dqPE5, dfdq_upd_prev_vec_out_AZ_dqPE5, dfdq_upd_prev_vec_out_LX_dqPE5, dfdq_upd_prev_vec_out_LY_dqPE5, dfdq_upd_prev_vec_out_LZ_dqPE5, dfdq_upd_prev_vec_out_AX_dqPE6, dfdq_upd_prev_vec_out_AY_dqPE6, dfdq_upd_prev_vec_out_AZ_dqPE6, dfdq_upd_prev_vec_out_LX_dqPE6, dfdq_upd_prev_vec_out_LY_dqPE6, dfdq_upd_prev_vec_out_LZ_dqPE6, dfdq_upd_prev_vec_out_AX_dqPE7, dfdq_upd_prev_vec_out_AY_dqPE7, dfdq_upd_prev_vec_out_AZ_dqPE7, dfdq_upd_prev_vec_out_LX_dqPE7, dfdq_upd_prev_vec_out_LY_dqPE7, dfdq_upd_prev_vec_out_LZ_dqPE7, dfdqd_upd_prev_vec_out_AX_dqdPE1, dfdqd_upd_prev_vec_out_AY_dqdPE1, dfdqd_upd_prev_vec_out_AZ_dqdPE1, dfdqd_upd_prev_vec_out_LX_dqdPE1, dfdqd_upd_prev_vec_out_LY_dqdPE1, dfdqd_upd_prev_vec_out_LZ_dqdPE1, dfdqd_upd_prev_vec_out_AX_dqdPE2, dfdqd_upd_prev_vec_out_AY_dqdPE2, dfdqd_upd_prev_vec_out_AZ_dqdPE2, dfdqd_upd_prev_vec_out_LX_dqdPE2, dfdqd_upd_prev_vec_out_LY_dqdPE2, dfdqd_upd_prev_vec_out_LZ_dqdPE2, dfdqd_upd_prev_vec_out_AX_dqdPE3, dfdqd_upd_prev_vec_out_AY_dqdPE3, dfdqd_upd_prev_vec_out_AZ_dqdPE3, dfdqd_upd_prev_vec_out_LX_dqdPE3, dfdqd_upd_prev_vec_out_LY_dqdPE3, dfdqd_upd_prev_vec_out_LZ_dqdPE3, dfdqd_upd_prev_vec_out_AX_dqdPE4, dfdqd_upd_prev_vec_out_AY_dqdPE4, dfdqd_upd_prev_vec_out_AZ_dqdPE4, dfdqd_upd_prev_vec_out_LX_dqdPE4, dfdqd_upd_prev_vec_out_LY_dqdPE4, dfdqd_upd_prev_vec_out_LZ_dqdPE4, dfdqd_upd_prev_vec_out_AX_dqdPE5, dfdqd_upd_prev_vec_out_AY_dqdPE5, dfdqd_upd_prev_vec_out_AZ_dqdPE5, dfdqd_upd_prev_vec_out_LX_dqdPE5, dfdqd_upd_prev_vec_out_LY_dqdPE5, dfdqd_upd_prev_vec_out_LZ_dqdPE5, dfdqd_upd_prev_vec_out_AX_dqdPE6, dfdqd_upd_prev_vec_out_AY_dqdPE6, dfdqd_upd_prev_vec_out_AZ_dqdPE6, dfdqd_upd_prev_vec_out_LX_dqdPE6, dfdqd_upd_prev_vec_out_LY_dqdPE6, dfdqd_upd_prev_vec_out_LZ_dqdPE6, dfdqd_upd_prev_vec_out_AX_dqdPE7, dfdqd_upd_prev_vec_out_AY_dqdPE7, dfdqd_upd_prev_vec_out_AZ_dqdPE7, dfdqd_upd_prev_vec_out_LX_dqdPE7, dfdqd_upd_prev_vec_out_LY_dqdPE7, dfdqd_upd_prev_vec_out_LZ_dqdPE7,
        minv_vec_out_R1_dqdPE1, minv_vec_out_R2_dqdPE1, minv_vec_out_R3_dqdPE1, minv_vec_out_R4_dqdPE1, minv_vec_out_R5_dqdPE1, minv_vec_out_R6_dqdPE1, minv_vec_out_R7_dqdPE1, minv_vec_out_R1_dqdPE2, minv_vec_out_R2_dqdPE2, minv_vec_out_R3_dqdPE2, minv_vec_out_R4_dqdPE2, minv_vec_out_R5_dqdPE2, minv_vec_out_R6_dqdPE2, minv_vec_out_R7_dqdPE2, minv_vec_out_R1_dqdPE3, minv_vec_out_R2_dqdPE3, minv_vec_out_R3_dqdPE3, minv_vec_out_R4_dqdPE3, minv_vec_out_R5_dqdPE3, minv_vec_out_R6_dqdPE3, minv_vec_out_R7_dqdPE3, minv_vec_out_R1_dqdPE4, minv_vec_out_R2_dqdPE4, minv_vec_out_R3_dqdPE4, minv_vec_out_R4_dqdPE4, minv_vec_out_R5_dqdPE4, minv_vec_out_R6_dqdPE4, minv_vec_out_R7_dqdPE4, minv_vec_out_R1_dqdPE5, minv_vec_out_R2_dqdPE5, minv_vec_out_R3_dqdPE5, minv_vec_out_R4_dqdPE5, minv_vec_out_R5_dqdPE5, minv_vec_out_R6_dqdPE5, minv_vec_out_R7_dqdPE5, minv_vec_out_R1_dqdPE6, minv_vec_out_R2_dqdPE6, minv_vec_out_R3_dqdPE6, minv_vec_out_R4_dqdPE6, minv_vec_out_R5_dqdPE6, minv_vec_out_R6_dqdPE6, minv_vec_out_R7_dqdPE6, minv_vec_out_R1_dqdPE7, minv_vec_out_R2_dqdPE7, minv_vec_out_R3_dqdPE7, minv_vec_out_R4_dqdPE7, minv_vec_out_R5_dqdPE7, minv_vec_out_R6_dqdPE7, minv_vec_out_R7_dqdPE7
    );

endmodule
