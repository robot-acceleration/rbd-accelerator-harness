result_vec[0] = new_minv_dtaudq[0][0];
result_vec[49+0] = new_minv_dtaudqd[0][0];
result_vec[1] = new_minv_dtaudq[0][1];
result_vec[49+1] = new_minv_dtaudqd[0][1];
result_vec[2] = new_minv_dtaudq[0][2];
result_vec[49+2] = new_minv_dtaudqd[0][2];
result_vec[3] = new_minv_dtaudq[0][3];
result_vec[49+3] = new_minv_dtaudqd[0][3];
result_vec[4] = new_minv_dtaudq[0][4];
result_vec[49+4] = new_minv_dtaudqd[0][4];
result_vec[5] = new_minv_dtaudq[0][5];
result_vec[49+5] = new_minv_dtaudqd[0][5];
result_vec[6] = new_minv_dtaudq[0][6];
result_vec[49+6] = new_minv_dtaudqd[0][6];
result_vec[7] = new_minv_dtaudq[1][0];
result_vec[49+7] = new_minv_dtaudqd[1][0];
result_vec[8] = new_minv_dtaudq[1][1];
result_vec[49+8] = new_minv_dtaudqd[1][1];
result_vec[9] = new_minv_dtaudq[1][2];
result_vec[49+9] = new_minv_dtaudqd[1][2];
result_vec[10] = new_minv_dtaudq[1][3];
result_vec[49+10] = new_minv_dtaudqd[1][3];
result_vec[11] = new_minv_dtaudq[1][4];
result_vec[49+11] = new_minv_dtaudqd[1][4];
result_vec[12] = new_minv_dtaudq[1][5];
result_vec[49+12] = new_minv_dtaudqd[1][5];
result_vec[13] = new_minv_dtaudq[1][6];
result_vec[49+13] = new_minv_dtaudqd[1][6];
result_vec[14] = new_minv_dtaudq[2][0];
result_vec[49+14] = new_minv_dtaudqd[2][0];
result_vec[15] = new_minv_dtaudq[2][1];
result_vec[49+15] = new_minv_dtaudqd[2][1];
result_vec[16] = new_minv_dtaudq[2][2];
result_vec[49+16] = new_minv_dtaudqd[2][2];
result_vec[17] = new_minv_dtaudq[2][3];
result_vec[49+17] = new_minv_dtaudqd[2][3];
result_vec[18] = new_minv_dtaudq[2][4];
result_vec[49+18] = new_minv_dtaudqd[2][4];
result_vec[19] = new_minv_dtaudq[2][5];
result_vec[49+19] = new_minv_dtaudqd[2][5];
result_vec[20] = new_minv_dtaudq[2][6];
result_vec[49+20] = new_minv_dtaudqd[2][6];
result_vec[21] = new_minv_dtaudq[3][0];
result_vec[49+21] = new_minv_dtaudqd[3][0];
result_vec[22] = new_minv_dtaudq[3][1];
result_vec[49+22] = new_minv_dtaudqd[3][1];
result_vec[23] = new_minv_dtaudq[3][2];
result_vec[49+23] = new_minv_dtaudqd[3][2];
result_vec[24] = new_minv_dtaudq[3][3];
result_vec[49+24] = new_minv_dtaudqd[3][3];
result_vec[25] = new_minv_dtaudq[3][4];
result_vec[49+25] = new_minv_dtaudqd[3][4];
result_vec[26] = new_minv_dtaudq[3][5];
result_vec[49+26] = new_minv_dtaudqd[3][5];
result_vec[27] = new_minv_dtaudq[3][6];
result_vec[49+27] = new_minv_dtaudqd[3][6];
result_vec[28] = new_minv_dtaudq[4][0];
result_vec[49+28] = new_minv_dtaudqd[4][0];
result_vec[29] = new_minv_dtaudq[4][1];
result_vec[49+29] = new_minv_dtaudqd[4][1];
result_vec[30] = new_minv_dtaudq[4][2];
result_vec[49+30] = new_minv_dtaudqd[4][2];
result_vec[31] = new_minv_dtaudq[4][3];
result_vec[49+31] = new_minv_dtaudqd[4][3];
result_vec[32] = new_minv_dtaudq[4][4];
result_vec[49+32] = new_minv_dtaudqd[4][4];
result_vec[33] = new_minv_dtaudq[4][5];
result_vec[49+33] = new_minv_dtaudqd[4][5];
result_vec[34] = new_minv_dtaudq[4][6];
result_vec[49+34] = new_minv_dtaudqd[4][6];
result_vec[35] = new_minv_dtaudq[5][0];
result_vec[49+35] = new_minv_dtaudqd[5][0];
result_vec[36] = new_minv_dtaudq[5][1];
result_vec[49+36] = new_minv_dtaudqd[5][1];
result_vec[37] = new_minv_dtaudq[5][2];
result_vec[49+37] = new_minv_dtaudqd[5][2];
result_vec[38] = new_minv_dtaudq[5][3];
result_vec[49+38] = new_minv_dtaudqd[5][3];
result_vec[39] = new_minv_dtaudq[5][4];
result_vec[49+39] = new_minv_dtaudqd[5][4];
result_vec[40] = new_minv_dtaudq[5][5];
result_vec[49+40] = new_minv_dtaudqd[5][5];
result_vec[41] = new_minv_dtaudq[5][6];
result_vec[49+41] = new_minv_dtaudqd[5][6];
result_vec[42] = new_minv_dtaudq[6][0];
result_vec[49+42] = new_minv_dtaudqd[6][0];
result_vec[43] = new_minv_dtaudq[6][1];
result_vec[49+43] = new_minv_dtaudqd[6][1];
result_vec[44] = new_minv_dtaudq[6][2];
result_vec[49+44] = new_minv_dtaudqd[6][2];
result_vec[45] = new_minv_dtaudq[6][3];
result_vec[49+45] = new_minv_dtaudqd[6][3];
result_vec[46] = new_minv_dtaudq[6][4];
result_vec[49+46] = new_minv_dtaudqd[6][4];
result_vec[47] = new_minv_dtaudq[6][5];
result_vec[49+47] = new_minv_dtaudqd[6][5];
result_vec[48] = new_minv_dtaudq[6][6];
result_vec[49+48] = new_minv_dtaudqd[6][6];
