// prevs for each PE
if (link_out_curr_PE != 0) begin
    dvda_prev[i] <= dvda_PE;
end
