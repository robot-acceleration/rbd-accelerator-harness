new_minv[0][0] = sparse_minv[0];
new_minv[0][1] = sparse_minv[1];
new_minv[0][2] = sparse_minv[2];
new_minv[0][3] = sparse_minv[3];
new_minv[0][4] = sparse_minv[4];
new_minv[0][5] = sparse_minv[5];
new_minv[0][6] = sparse_minv[6];
new_minv[1][0] = sparse_minv[7];
new_minv[1][1] = sparse_minv[8];
new_minv[1][2] = sparse_minv[9];
new_minv[1][3] = sparse_minv[10];
new_minv[1][4] = sparse_minv[11];
new_minv[1][5] = sparse_minv[12];
new_minv[1][6] = sparse_minv[13];
new_minv[2][0] = sparse_minv[14];
new_minv[2][1] = sparse_minv[15];
new_minv[2][2] = sparse_minv[16];
new_minv[2][3] = sparse_minv[17];
new_minv[2][4] = sparse_minv[18];
new_minv[2][5] = sparse_minv[19];
new_minv[2][6] = sparse_minv[20];
new_minv[3][0] = sparse_minv[21];
new_minv[3][1] = sparse_minv[22];
new_minv[3][2] = sparse_minv[23];
new_minv[3][3] = sparse_minv[24];
new_minv[3][4] = sparse_minv[25];
new_minv[3][5] = sparse_minv[26];
new_minv[3][6] = sparse_minv[27];
new_minv[4][0] = sparse_minv[28];
new_minv[4][1] = sparse_minv[29];
new_minv[4][2] = sparse_minv[30];
new_minv[4][3] = sparse_minv[31];
new_minv[4][4] = sparse_minv[32];
new_minv[4][5] = sparse_minv[33];
new_minv[4][6] = sparse_minv[34];
new_minv[5][0] = sparse_minv[35];
new_minv[5][1] = sparse_minv[36];
new_minv[5][2] = sparse_minv[37];
new_minv[5][3] = sparse_minv[38];
new_minv[5][4] = sparse_minv[39];
new_minv[5][5] = sparse_minv[40];
new_minv[5][6] = sparse_minv[41];
new_minv[6][0] = sparse_minv[42];
new_minv[6][1] = sparse_minv[43];
new_minv[6][2] = sparse_minv[44];
new_minv[6][3] = sparse_minv[45];
new_minv[6][4] = sparse_minv[46];
new_minv[6][5] = sparse_minv[47];
new_minv[6][6] = sparse_minv[48];
